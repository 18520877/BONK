// Convolution Kernel 3x3, Stride = 2, Padding = 0. 
//Input = 299x299x3, Output = 147x147x96.

module Conv2d_1a_3x3_32
#(parameter D = 220,
  parameter DATA_WIDTH = 32)
(
     //input
    	input clk,
    	input reset,
    	input valid_in_1, valid_in_2, valid_in_3,
    	input [DATA_WIDTH-1:0] pxl_in_1, pxl_in_2, pxl_in_3,
    
output [DATA_WIDTH-1:0] pxl_out_1 , pxl_out_2 , pxl_out_3 , pxl_out_4 , pxl_out_5 , pxl_out_6 , pxl_out_7 , pxl_out_8 , pxl_out_9 , pxl_out_10,
                        pxl_out_11, pxl_out_12, pxl_out_13, pxl_out_14, pxl_out_15, pxl_out_16, pxl_out_17, pxl_out_18, pxl_out_19, pxl_out_20,
	                      pxl_out_21, pxl_out_22, pxl_out_23, pxl_out_24, pxl_out_25, pxl_out_26, pxl_out_27, pxl_out_28, pxl_out_29, pxl_out_30,
                        pxl_out_31, pxl_out_32, pxl_out_33, pxl_out_34, pxl_out_35, pxl_out_36, pxl_out_37, pxl_out_38, pxl_out_39, pxl_out_40,
                        pxl_out_41, pxl_out_42, pxl_out_43, pxl_out_44, pxl_out_45, pxl_out_46, pxl_out_47, pxl_out_48, pxl_out_49, pxl_out_50,
                        pxl_out_51, pxl_out_52, pxl_out_53, pxl_out_54, pxl_out_55, pxl_out_56, pxl_out_57, pxl_out_58, pxl_out_59, pxl_out_60,
                        pxl_out_61, pxl_out_62, pxl_out_63, pxl_out_64, pxl_out_65, pxl_out_66, pxl_out_67, pxl_out_68, pxl_out_69, pxl_out_70,
                        pxl_out_71, pxl_out_72, pxl_out_73, pxl_out_74, pxl_out_75, pxl_out_76, pxl_out_77, pxl_out_78, pxl_out_79, pxl_out_80,
                        pxl_out_81, pxl_out_82, pxl_out_83, pxl_out_84, pxl_out_85, pxl_out_86, pxl_out_87, pxl_out_88, pxl_out_89, pxl_out_90,
                        pxl_out_91, pxl_out_92, pxl_out_93, pxl_out_94, pxl_out_95, pxl_out_96,   
                                              
	               output valid_out_1 , valid_out_2 , valid_out_3 , valid_out_4 , valid_out_5 , valid_out_6 , valid_out_7 , valid_out_8 , valid_out_9 , valid_out_10,
                        valid_out_11, valid_out_12, valid_out_13, valid_out_14, valid_out_15, valid_out_16, valid_out_17, valid_out_18, valid_out_19, valid_out_20,
	                      valid_out_21, valid_out_22, valid_out_23, valid_out_24, valid_out_25, valid_out_26, valid_out_27, valid_out_28, valid_out_29, valid_out_30,
                        valid_out_31, valid_out_32, valid_out_33, valid_out_34, valid_out_35, valid_out_36, valid_out_37, valid_out_38, valid_out_39, valid_out_40,
                        valid_out_41, valid_out_42, valid_out_43, valid_out_44, valid_out_45, valid_out_46, valid_out_47, valid_out_48, valid_out_49, valid_out_50,
                        valid_out_51, valid_out_52, valid_out_53, valid_out_54, valid_out_55, valid_out_56, valid_out_57, valid_out_58, valid_out_59, valid_out_60,
                        valid_out_61, valid_out_62, valid_out_63, valid_out_64, valid_out_65, valid_out_66, valid_out_67, valid_out_68, valid_out_69, valid_out_70,
                        valid_out_71, valid_out_72, valid_out_73, valid_out_74, valid_out_75, valid_out_76, valid_out_77, valid_out_78, valid_out_79, valid_out_80,
                        valid_out_81, valid_out_82, valid_out_83, valid_out_84, valid_out_85, valid_out_86, valid_out_87, valid_out_88, valid_out_89, valid_out_90,
                        valid_out_91, valid_out_92, valid_out_93, valid_out_94, valid_out_95, valid_out_96  
	     
);

//Channel 1
conv_33_s2 #(D, DATA_WIDTH) x1(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b10111110001001110100011100001000),
.kernel_01(32'b10111011110010100011010100101100),
.kernel_02(32'b00111110000001100010111110100011),
.kernel_03(32'b00111101000101110111011100111000),
.kernel_04(32'b10111110000000000110011001011010),
.kernel_05(32'b00111101011001110110001110100000),
.kernel_06(32'b10111101000010001110001100001111),
.kernel_07(32'b00111101000111011011100110101011),
.kernel_08(32'b10111110000100011011101100110111),
.pxl_out(pxl_out_1), .valid_out(valid_out_1) );

//Channel 2
conv_33_s2 #(D, DATA_WIDTH) x2(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b10111110111011100111011111001010),
.kernel_01(32'b00111100111011000111011110111110),
.kernel_02(32'b10111110011010110111100010011001),
.kernel_03(32'b00111110100101100101111001101111),
.kernel_04(32'b00111110101111010111010110100000),
.kernel_05(32'b00111100001010111100111011111010),
.kernel_06(32'b10111101011100111110111111010000),
.kernel_07(32'b00111011100000111111000001000011),
.kernel_08(32'b10111111001010001011111000101101),
.pxl_out(pxl_out_2), .valid_out(valid_out_2) );

//Channel 3
conv_33_s2 #(D, DATA_WIDTH) x3(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b00111110111101001100011110110000),
.kernel_01(32'b00111110100000100110101110101010),
.kernel_02(32'b10111011101011110100101001111110),
.kernel_03(32'b00111110111101111001100111000001),
.kernel_04(32'b10111110010101100011010110110111),
.kernel_05(32'b00111111000101001100001100000000),
.kernel_06(32'b10111100010111011000001000000110),
.kernel_07(32'b00111110110111011010001111010011),
.kernel_08(32'b10111110110100010100101101111000),
.pxl_out(pxl_out_3), .valid_out(valid_out_3) );

//Channel 4
conv_33_s2 #(D, DATA_WIDTH) x4(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b00111110000001000110110000110010),
.kernel_01(32'b00111110100101011011111101110100),
.kernel_02(32'b00111110000001001111110011010100),
.kernel_03(32'b10111101100011111000011011001101),
.kernel_04(32'b10111110010000010110001110111111),
.kernel_05(32'b00111100100100000111111010110001),
.kernel_06(32'b00111100100100111110011101101110),
.kernel_07(32'b10111101011110000111100000011110),
.kernel_08(32'b00111110000101001111100011100000),
.pxl_out(pxl_out_4), .valid_out(valid_out_4) );

//Channel 5
conv_33_s2 #(D, DATA_WIDTH) x5(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b10111101011110001100111011000101),
.kernel_01(32'b00111100111010001000011110011111),
.kernel_02(32'b10111101001101110100010011001001),
.kernel_03(32'b10111101010001010100001100011100),
.kernel_04(32'b00111101001111101011110000010111),
.kernel_05(32'b10111111000110011101000011111011),
.kernel_06(32'b10111101001100110100000010100100),
.kernel_07(32'b00111111000010101110001111101101),
.kernel_08(32'b00111110110101110110100011010100),
.pxl_out(pxl_out_5), .valid_out(valid_out_5) );

//Channel 6
conv_33_s2 #(D, DATA_WIDTH) x6(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b00111110111010011110010011010001),
.kernel_01(32'b10111101010001011101101100010111),
.kernel_02(32'b00111101111111000000010101010000),
.kernel_03(32'b10111110101111000100011000110101),
.kernel_04(32'b10111111000110001101001000011010),
.kernel_05(32'b10111110110000111111101110001110),
.kernel_06(32'b10111110001011010001111010001001),
.kernel_07(32'b00111101001000110111000011000111),
.kernel_08(32'b00111111000000100000000000110100),
.pxl_out(pxl_out_6), .valid_out(valid_out_6) );

//Channel 7
conv_33_s2 #(D, DATA_WIDTH) x7(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b00111100100110001001111001100000),
.kernel_01(32'b00111111001101010111100111010010),
.kernel_02(32'b00111000011100111010100111001100),
.kernel_03(32'b00111011110111001010101110011011),
.kernel_04(32'b10111110110011100010001111000111),
.kernel_05(32'b00111110000001010111101001111010),
.kernel_06(32'b00111110011011011001001100000110),
.kernel_07(32'b00111110011111111110111100110111),
.kernel_08(32'b10111100110001011100010011010011),
.pxl_out(pxl_out_7), .valid_out(valid_out_7) );

//Channel 8
conv_33_s2 #(D, DATA_WIDTH) x8(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b00111110001110011100010110011111),
.kernel_01(32'b00111011110010111110101011000101),
.kernel_02(32'b00111101100010010001101111000110),
.kernel_03(32'b10111101001000001110010011011000),
.kernel_04(32'b00111110001011000101011001101011),
.kernel_05(32'b00111101000110101010011110010011),
.kernel_06(32'b10111101101011011010110110101111),
.kernel_07(32'b00111101101100111111100110110110),
.kernel_08(32'b10111110011111100111010110001010),
.pxl_out(pxl_out_8), .valid_out(valid_out_8) );

//Channel 9
conv_33_s2 #(D, DATA_WIDTH) x9(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b00111110000111010001001110101101),
.kernel_01(32'b10111110100011011011110110001110),
.kernel_02(32'b10111110011111001101100101010100),
.kernel_03(32'b10111110100101110110011101101000),
.kernel_04(32'b00111110001111100000001100000010),
.kernel_05(32'b00111101110111111111000000100001),
.kernel_06(32'b00111100000110000001111011100111),
.kernel_07(32'b10111101011111100001010001100101),
.kernel_08(32'b00111110101100100111110010101110),
.pxl_out(pxl_out_9), .valid_out(valid_out_9) );

//Channel 10
conv_33_s2 #(D, DATA_WIDTH) x10(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b10111110100110101100000110101110),
.kernel_01(32'b10111101101001110100001010000111),
.kernel_02(32'b10111101111100111011001000110011),
.kernel_03(32'b10111101111000101010111010001010),
.kernel_04(32'b00111110101010110100101010111001),
.kernel_05(32'b00111110000011100011011111110101),
.kernel_06(32'b00111110011101101011011100010010),
.kernel_07(32'b10111101100010011111000001101001),
.kernel_08(32'b10111110101011001001011101000110),
.pxl_out(pxl_out_10), .valid_out(valid_out_10) );

//Channel 11
conv_33_s2 #(D, DATA_WIDTH) x11(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b10111110110010111110101010001000),
.kernel_01(32'b10111110101000000111111010001111),
.kernel_02(32'b00111101100001001000001001000111),
.kernel_03(32'b00111110100011100001110100011011),
.kernel_04(32'b10111101100001000101110110100001),
.kernel_05(32'b00111101101000101110101100111111),
.kernel_06(32'b10111111000100001001100001001000),
.kernel_07(32'b10111101000100111001001001100010),
.kernel_08(32'b00111110100000001111110100110111),
.pxl_out(pxl_out_11), .valid_out(valid_out_11) );

//Channel 12
conv_33_s2 #(D, DATA_WIDTH) x12(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b00111101101111011000110001111001),
.kernel_01(32'b00111101100110010110010111100010),
.kernel_02(32'b10111101010110000111100101101001),
.kernel_03(32'b00111110001000010011111101101011),
.kernel_04(32'b10111101001010101100011101111101),
.kernel_05(32'b10111110011110011011101001010101),
.kernel_06(32'b10111111100001000111100000011110),
.kernel_07(32'b10111100000000001110011000111111),
.kernel_08(32'b10111110100000001101100111101100),
.pxl_out(pxl_out_12), .valid_out(valid_out_12) );

//Channel 13
conv_33_s2 #(D, DATA_WIDTH) x13(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b00111101010011011011001010110101),
.kernel_01(32'b00111111010111001011100000110111),
.kernel_02(32'b00111101111010000111010101001111),
.kernel_03(32'b10111101110100100011010011100000),
.kernel_04(32'b00111101000111101111011000001101),
.kernel_05(32'b00111111000101010110011100011100),
.kernel_06(32'b00111111001000011101111001110001),
.kernel_07(32'b00111110100001011110100111101000),
.kernel_08(32'b00111100110011101011101100001110),
.pxl_out(pxl_out_13), .valid_out(valid_out_13) );

//Channel 14
conv_33_s2 #(D, DATA_WIDTH) x14(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b00111111011110111011010010011011),
.kernel_01(32'b10111110100100110101011101111101),
.kernel_02(32'b00111101011110100011101010100100),
.kernel_03(32'b00111100010001000011100110001000),
.kernel_04(32'b00111111001001011100011100010111),
.kernel_05(32'b10111110100001010110011010110011),
.kernel_06(32'b00111110101010011001011111011001),
.kernel_07(32'b10111111000101011101111001100001),
.kernel_08(32'b10111110101000100000111000001001),
.pxl_out(pxl_out_14), .valid_out(valid_out_14) );

//Channel 15
conv_33_s2 #(D, DATA_WIDTH) x15(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b00111110100000001000010110010000),
.kernel_01(32'b10111110110001111001111011001010),
.kernel_02(32'b00111101100000111011110001100101),
.kernel_03(32'b00111100111010100100111111001100),
.kernel_04(32'b00111011101000010001001111010100),
.kernel_05(32'b00111101100100111011100100110000),
.kernel_06(32'b00111101101010111101100011100000),
.kernel_07(32'b10111101011100000001111110000001),
.kernel_08(32'b00111101110011000000100111111000),
.pxl_out(pxl_out_15), .valid_out(valid_out_15) );

//Channel 16
conv_33_s2 #(D, DATA_WIDTH) x16(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b10111101110000100100101110110101),
.kernel_01(32'b00111101010110011100111001110101),
.kernel_02(32'b10111111101001111111101101111000),
.kernel_03(32'b00111110000110100100000000111111),
.kernel_04(32'b00111111010101011000101011000111),
.kernel_05(32'b00111101010100011110101001100010),
.kernel_06(32'b00111111100110001111110111111011),
.kernel_07(32'b10111101110000111100100100110110),
.kernel_08(32'b00111110010110011000011100010000),
.pxl_out(pxl_out_16), .valid_out(valid_out_16) );

//Channel 17
conv_33_s2 #(D, DATA_WIDTH) x17(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b10111111000101100111110010111010),
.kernel_01(32'b00111110111111111111000101000101),
.kernel_02(32'b10111111000110011010011101000101),
.kernel_03(32'b10111110001011010110001010111110),
.kernel_04(32'b10111100110001001001100111110001),
.kernel_05(32'b00111111100010011100001100001100),
.kernel_06(32'b00111100000010110110011011011000),
.kernel_07(32'b00111101101001010010110111001010),
.kernel_08(32'b00111100110001100100110111010000),
.pxl_out(pxl_out_17), .valid_out(valid_out_17) );

//Channel 18
conv_33_s2 #(D, DATA_WIDTH) x18(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b10111110000000011000110111001101),
.kernel_01(32'b10111110000100000001011101000101),
.kernel_02(32'b00111110100011100001011100001101),
.kernel_03(32'b10111111000111001000010101111010),
.kernel_04(32'b10111110011010111110111110100000),
.kernel_05(32'b00111110100010001000011011000000),
.kernel_06(32'b00111110100011001111000010001000),
.kernel_07(32'b00111100101011100000110111110110),
.kernel_08(32'b00111101000010111001100010100101),
.pxl_out(pxl_out_18), .valid_out(valid_out_18) );

//Channel 19
conv_33_s2 #(D, DATA_WIDTH) x19(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b00111101000101011000000110010000),
.kernel_01(32'b00111101111011111001111111110011),
.kernel_02(32'b00111101010100000101001101100101),
.kernel_03(32'b10111101101110010101110000000001),
.kernel_04(32'b00111110000010111000101010101110),
.kernel_05(32'b10111110110101101100100000111101),
.kernel_06(32'b00111101111111000101101111101001),
.kernel_07(32'b10111111001011110100111110000100),
.kernel_08(32'b10111011100011101100110010001001),
.pxl_out(pxl_out_19), .valid_out(valid_out_19) );

//Channel 20
conv_33_s2 #(D, DATA_WIDTH) x20(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b10111111000011001101100101111010),
.kernel_01(32'b00111101010100011011010011011110),
.kernel_02(32'b00111111001000000011010011010010),
.kernel_03(32'b10111101000011110001001010101110),
.kernel_04(32'b10111101100101001111111111010110),
.kernel_05(32'b00111111000100011001111100001100),
.kernel_06(32'b00111110100110011010000001100101),
.kernel_07(32'b10111101101011001111001101000001),
.kernel_08(32'b10111101100010001100101000101000),
.pxl_out(pxl_out_20), .valid_out(valid_out_20) );

//Channel 21
conv_33_s2 #(D, DATA_WIDTH) x21(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b10111110100010001000001111011100),
.kernel_01(32'b00111111010010000000111011100100),
.kernel_02(32'b00111110101001111010111010011000),
.kernel_03(32'b00111101000110001110001101001001),
.kernel_04(32'b10111110000000110001010000001110),
.kernel_05(32'b10111111000100010101000100001011),
.kernel_06(32'b10111110010100110001000010010001),
.kernel_07(32'b10111110111011110101010111100001),
.kernel_08(32'b10111110101111110100101101100101),
.pxl_out(pxl_out_21), .valid_out(valid_out_21) );

//Channel 22
conv_33_s2 #(D, DATA_WIDTH) x22(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b10111110100001001000001111111101),
.kernel_01(32'b00111110001010101111100001101011),
.kernel_02(32'b00111110000111100101001100101010),
.kernel_03(32'b10111101001011001111011101101100),
.kernel_04(32'b10111101100100111000111101000011),
.kernel_05(32'b00111110000011110000000010010000),
.kernel_06(32'b00111100110100010101100101111111),
.kernel_07(32'b00111101011010000000110011100000),
.kernel_08(32'b00111101010101011111010101100011),
.pxl_out(pxl_out_22), .valid_out(valid_out_22) );

//Channel 23
conv_33_s2 #(D, DATA_WIDTH) x23(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b00111110000101101110110111010000),
.kernel_01(32'b10111100101001100011010101000011),
.kernel_02(32'b10111101101001100010001110011111),
.kernel_03(32'b10111111000001101101100110000000),
.kernel_04(32'b10111110011011000001000001110000),
.kernel_05(32'b10111101111010011111000100101101),
.kernel_06(32'b10111110101011001000100010011101),
.kernel_07(32'b00111111000001001100011010011011),
.kernel_08(32'b10111100000101111101110111101111),
.pxl_out(pxl_out_23), .valid_out(valid_out_23) );

//Channel 24
conv_33_s2 #(D, DATA_WIDTH) x24(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b00111100110100010110101111010101),
.kernel_01(32'b00111101100011100011001001110001),
.kernel_02(32'b00111101000011000010010011110011),
.kernel_03(32'b00111110100101001101111000100010),
.kernel_04(32'b00111110001110100010101100110111),
.kernel_05(32'b10111100010000111111110011110110),
.kernel_06(32'b00111110111110011001111001010111),
.kernel_07(32'b10111110011111011011100000000110),
.kernel_08(32'b10111111001000000100100101001011),
.pxl_out(pxl_out_24), .valid_out(valid_out_24) );

//Channel 25
conv_33_s2 #(D, DATA_WIDTH) x25(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b00111100000111001110010000111001),
.kernel_01(32'b00111110101001101100001110101001),
.kernel_02(32'b00111110101100000110100101001110),
.kernel_03(32'b00111110001001011101110000110011),
.kernel_04(32'b00111110110101011010111111100100),
.kernel_05(32'b10111110101101000011011011001100),
.kernel_06(32'b10111110100000111011100100110000),
.kernel_07(32'b10111101010010010101111101010100),
.kernel_08(32'b10111101010010100000110100101010),
.pxl_out(pxl_out_25), .valid_out(valid_out_25) );

//Channel 26
conv_33_s2 #(D, DATA_WIDTH) x26(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b00111100101100101110111000011101),
.kernel_01(32'b00111101001001000010100100011011),
.kernel_02(32'b00111011100111101111001001010011),
.kernel_03(32'b10111010100000111100101000110000),
.kernel_04(32'b00111100110101000111010101101001),
.kernel_05(32'b00111101011010010110111111010111),
.kernel_06(32'b10111101100111011100001111101111),
.kernel_07(32'b00111101110100100001000100101010),
.kernel_08(32'b10111111001000101001101111000010),
.pxl_out(pxl_out_26), .valid_out(valid_out_26) );

//Channel 27
conv_33_s2 #(D, DATA_WIDTH) x27(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b00111110010000101101101000000001),
.kernel_01(32'b00111110111101000111010011000110),
.kernel_02(32'b10111110110111101011011010111001),
.kernel_03(32'b00111111001101001101110111101010),
.kernel_04(32'b10111101100000000011101010110001),
.kernel_05(32'b00111101100011111101000100111111),
.kernel_06(32'b10111110110011111110000111001010),
.kernel_07(32'b00111101110110111010100000010110),
.kernel_08(32'b10111110101000101110001010010000),
.pxl_out(pxl_out_27), .valid_out(valid_out_27) );

//Channel 28
conv_33_s2 #(D, DATA_WIDTH) x28(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b10111110001011010101101101001100),
.kernel_01(32'b00111101001011000100111001101001),
.kernel_02(32'b00111111000010111101000111110001),
.kernel_03(32'b00111101001001001010001101011011),
.kernel_04(32'b10111111010001010000101100011100),
.kernel_05(32'b10111011000001010101100111011000),
.kernel_06(32'b10111101100000001100111111000100),
.kernel_07(32'b00111110110011101111111010000001),
.kernel_08(32'b00111110000100111000001011011001),
.pxl_out(pxl_out_28), .valid_out(valid_out_28) );

//Channel 29
conv_33_s2 #(D, DATA_WIDTH) x29(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b00111110110001001100010100110000),
.kernel_01(32'b10111110101010101101010000111110),
.kernel_02(32'b10111110011000010010100010100101),
.kernel_03(32'b00111110000101011100001011101100),
.kernel_04(32'b00111011100000000111011001011001),
.kernel_05(32'b10111100001110110011010101000111),
.kernel_06(32'b00111100000001000100111100000011),
.kernel_07(32'b10111101101000010111100011100110),
.kernel_08(32'b10111101111100110010101111110101),
.pxl_out(pxl_out_29), .valid_out(valid_out_29) );

//Channel 30
conv_33_s2 #(D, DATA_WIDTH) x30(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b10111101100010101000101101111001),
.kernel_01(32'b00111101101011000001011110111101),
.kernel_02(32'b10111110011110101011010101001111),
.kernel_03(32'b00111110000101101100011110100100),
.kernel_04(32'b10111110101111010110101010010100),
.kernel_05(32'b00111110101010000000100100011001),
.kernel_06(32'b10111110110001101000110001100010),
.kernel_07(32'b10111110100001011001100101101110),
.kernel_08(32'b00111110101011000101011000111101),
.pxl_out(pxl_out_30), .valid_out(valid_out_30) );

//Channel 31
conv_33_s2 #(D, DATA_WIDTH) x31(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b00111100101000101000000110010010),
.kernel_01(32'b10111110000000101101000100101011),
.kernel_02(32'b00111110101010010010010110010000),
.kernel_03(32'b00111101100001101100101100000011),
.kernel_04(32'b00111100111100110011011111101101),
.kernel_05(32'b10111101110001110111011100100111),
.kernel_06(32'b10111101101010100000111100010010),
.kernel_07(32'b00111110101010000111011100111000),
.kernel_08(32'b00111110100011110100111100010011),
.pxl_out(pxl_out_31), .valid_out(valid_out_31) );

//Channel 32
conv_33_s2 #(D, DATA_WIDTH) x32(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b10111110100111000010000101010101),
.kernel_01(32'b10111101110110000000010010011101),
.kernel_02(32'b10111110101100000010000111001101),
.kernel_03(32'b00111110101011011100101001010100),
.kernel_04(32'b10111110001101001001111011111101),
.kernel_05(32'b00111110001100100001111011101001),
.kernel_06(32'b10111110110000000101010001000100),
.kernel_07(32'b10111110000000110000000100011110),
.kernel_08(32'b10111101000010001001011111100101),
.pxl_out(pxl_out_32), .valid_out(valid_out_32) );

//Channel 33
conv_33_s2 #(D, DATA_WIDTH) x33(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b00111110000111000110110100111010),
.kernel_01(32'b10111101101010000101100101111001),
.kernel_02(32'b00111110011110110001111101011111),
.kernel_03(32'b00111110001000001000101111000001),
.kernel_04(32'b10111111001110010010110011011110),
.kernel_05(32'b10111110111100011011100100100011),
.kernel_06(32'b10111110101100001001101100101011),
.kernel_07(32'b00111101101010011111110001100110),
.kernel_08(32'b10111110001011100011011010000100),
.pxl_out(pxl_out_33), .valid_out(valid_out_33) );

//Channel 34
conv_33_s2 #(D, DATA_WIDTH) x34(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b00111110000100001011100000001101),
.kernel_01(32'b00111110010110001000101010111010),
.kernel_02(32'b10111110100010101111001111111100),
.kernel_03(32'b00111110011011111111001111011001),
.kernel_04(32'b00111100111010011111101100110001),
.kernel_05(32'b00111110001100100010001000111101),
.kernel_06(32'b10111110100011010111110111001100),
.kernel_07(32'b00111101110010001011001010110000),
.kernel_08(32'b10111111011010000111110001101000),
.pxl_out(pxl_out_34), .valid_out(valid_out_34) );

//Channel 35
conv_33_s2 #(D, DATA_WIDTH) x35(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b00111111000100011000110101111111),
.kernel_01(32'b10111110000011000010010101101110),
.kernel_02(32'b10111101001101111111110110011001),
.kernel_03(32'b10111110111011110110110011001010),
.kernel_04(32'b10111110001001001101011010011011),
.kernel_05(32'b00111110110000101100100110001110),
.kernel_06(32'b00111111000010001011101010011011),
.kernel_07(32'b00111111001011010001011001110110),
.kernel_08(32'b10111111001100001010111101011010),
.pxl_out(pxl_out_35), .valid_out(valid_out_35) );

//Channel 36
conv_33_s2 #(D, DATA_WIDTH) x36(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b00111110110100000010101000111101),
.kernel_01(32'b00111111000011110111010110101001),
.kernel_02(32'b00111110111111100001111110010101),
.kernel_03(32'b00111110111000101110100110010011),
.kernel_04(32'b10111111000101111111001001110000),
.kernel_05(32'b10111101100011111010000100111111),
.kernel_06(32'b10111101000001001100010010110110),
.kernel_07(32'b10111101111110011110110101001010),
.kernel_08(32'b00111110001110101011100100010001),
.pxl_out(pxl_out_36), .valid_out(valid_out_36) );

//Channel 37
conv_33_s2 #(D, DATA_WIDTH) x37(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b10111111010101010010101001000111),
.kernel_01(32'b10111110111001111000101111111001),
.kernel_02(32'b10111110100010001110000110000001),
.kernel_03(32'b00111101011110110001101001000010),
.kernel_04(32'b10111100110001101110010000010101),
.kernel_05(32'b00111110000011000011000010000001),
.kernel_06(32'b00111110000111111111101101011000),
.kernel_07(32'b00111111010011011110001010111111),
.kernel_08(32'b00111110101000100110111111100111),
.pxl_out(pxl_out_37), .valid_out(valid_out_37) );

//Channel 38
conv_33_s2 #(D, DATA_WIDTH) x38(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b00111100110010000100100111011001),
.kernel_01(32'b10111101101110011001001000010110),
.kernel_02(32'b00111110100111001110001100111000),
.kernel_03(32'b10111111000110101000011100110011),
.kernel_04(32'b10111111010111011100100010110111),
.kernel_05(32'b10111111000000010110101101000000),
.kernel_06(32'b00111101001110101111100111001011),
.kernel_07(32'b10111100000111001001000010011010),
.kernel_08(32'b10111111000000110111110111101000),
.pxl_out(pxl_out_38), .valid_out(valid_out_38) );

//Channel 39
conv_33_s2 #(D, DATA_WIDTH) x39(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b00111101100000101000001000011101),
.kernel_01(32'b00111110111100011111100001001011),
.kernel_02(32'b00111110111011100011001001011111),
.kernel_03(32'b10111110010000101001000010000110),
.kernel_04(32'b10111111001010110001100100100101),
.kernel_05(32'b00111110100111111000111111000000),
.kernel_06(32'b00111111000111100110010010010011),
.kernel_07(32'b00111111001001100010101001011100),
.kernel_08(32'b00111111000001011100001011010100),
.pxl_out(pxl_out_39), .valid_out(valid_out_39) );

//Channel 40
conv_33_s2 #(D, DATA_WIDTH) x40(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b00111110101010100000110111100000),
.kernel_01(32'b10111101001001001010101101011101),
.kernel_02(32'b00111101110101100010101011000101),
.kernel_03(32'b10111100001110000111101110111000),
.kernel_04(32'b00111110011100011011110001110011),
.kernel_05(32'b10111110101100000101100000101001),
.kernel_06(32'b10111110011000010110110101101011),
.kernel_07(32'b10111100100000000111000011100110),
.kernel_08(32'b00111101000011011110011100010001),
.pxl_out(pxl_out_40), .valid_out(valid_out_40) );

//Channel 41
conv_33_s2 #(D, DATA_WIDTH) x41(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b00111101101110111100100001001010),
.kernel_01(32'b00111101100100011000100100000001),
.kernel_02(32'b10111110110010101011100011110111),
.kernel_03(32'b10111111000010110101011011001100),
.kernel_04(32'b00111110001000110010011000001110),
.kernel_05(32'b10111011000100101011000110010000),
.kernel_06(32'b10111101011001111000101011000100),
.kernel_07(32'b10111101110110101101111100111011),
.kernel_08(32'b00111110111111100001001001011111),
.pxl_out(pxl_out_41), .valid_out(valid_out_41) );

//Channel 42
conv_33_s2 #(D, DATA_WIDTH) x42(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b10111111000011111110100011001100),
.kernel_01(32'b10111101010011011000000111110111),
.kernel_02(32'b00111100011100110010101100000111),
.kernel_03(32'b10111110001011101000111111011010),
.kernel_04(32'b10111110100010100101101010100101),
.kernel_05(32'b00111110100101101100000111111101),
.kernel_06(32'b00111110001000111001110111011111),
.kernel_07(32'b00111110101101001000000100110100),
.kernel_08(32'b10111111001000100010011010101000),
.pxl_out(pxl_out_42), .valid_out(valid_out_42) );

//Channel 43
conv_33_s2 #(D, DATA_WIDTH) x43(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b10111111001010001011011000001010),
.kernel_01(32'b10111110111110110100011111001100),
.kernel_02(32'b00111110101111101001100010111100),
.kernel_03(32'b00111111000000010001011000001000),
.kernel_04(32'b00111110010000101000010110011110),
.kernel_05(32'b00111110100011100011101001100101),
.kernel_06(32'b10111101111100110110111000011000),
.kernel_07(32'b10111101110101010110111000100000),
.kernel_08(32'b00111110110100010111011100000110),
.pxl_out(pxl_out_43), .valid_out(valid_out_43) );

//Channel 44
conv_33_s2 #(D, DATA_WIDTH) x44(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b00111110000110110100001100010111),
.kernel_01(32'b00111100011000001000111000010111),
.kernel_02(32'b10111111011100110110110001000101),
.kernel_03(32'b00111101110110110010011011111010),
.kernel_04(32'b00111101110100001000011111111000),
.kernel_05(32'b10111110100000011100100010010101),
.kernel_06(32'b00111110101111001011100001110101),
.kernel_07(32'b00111101101111100001001111011011),
.kernel_08(32'b10111110110011001101101010100001),
.pxl_out(pxl_out_44), .valid_out(valid_out_44) );

//Channel 45
conv_33_s2 #(D, DATA_WIDTH) x45(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b00111101100111011100101001101011),
.kernel_01(32'b00111011010001001101111000101101),
.kernel_02(32'b00111110100011011001111100011001),
.kernel_03(32'b10111110110111010001011110110011),
.kernel_04(32'b00111110000011100000100010011110),
.kernel_05(32'b00111111011011101110011110100001),
.kernel_06(32'b00111111010001000110101001000001),
.kernel_07(32'b10111110111110100011101111011100),
.kernel_08(32'b10111101010011011011110110111101),
.pxl_out(pxl_out_45), .valid_out(valid_out_45) );

//Channel 46
conv_33_s2 #(D, DATA_WIDTH) x46(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b10111111011001110000010000111110),
.kernel_01(32'b10111110100010011010100110010001),
.kernel_02(32'b00111100110110011010011110001101),
.kernel_03(32'b00111111011001001110110111000000),
.kernel_04(32'b00111111100001101111111001010100),
.kernel_05(32'b10111110111001111001000001011100),
.kernel_06(32'b00111111001110101101011111001011),
.kernel_07(32'b10111111100111111001110101010101),
.kernel_08(32'b10111110111111000110110111111101),
.pxl_out(pxl_out_46), .valid_out(valid_out_46) );

//Channel 47
conv_33_s2 #(D, DATA_WIDTH) x47(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b00111111000011011101101001101000),
.kernel_01(32'b10111111011111000010111000101011),
.kernel_02(32'b10111100011110010111111000000111),
.kernel_03(32'b10111101110110100001101100110101),
.kernel_04(32'b10111101100001001101000100110110),
.kernel_05(32'b00111101100011100001000100110111),
.kernel_06(32'b00111100101000011100011010001000),
.kernel_07(32'b10111111011111100110010011110010),
.kernel_08(32'b00111101000111110101100111010101),
.pxl_out(pxl_out_47), .valid_out(valid_out_47) );

//Channel 48
conv_33_s2 #(D, DATA_WIDTH) x48(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b00111101000111011111001101001110),
.kernel_01(32'b10111101100111100111110101000001),
.kernel_02(32'b00111110101100101010111011001010),
.kernel_03(32'b00111110001101011101111000111011),
.kernel_04(32'b00111111100110111101100000011011),
.kernel_05(32'b00111101101011100100010110100111),
.kernel_06(32'b00111101001110101110101011011100),
.kernel_07(32'b10111101111111101100111110001001),
.kernel_08(32'b00111110111111110101101101101101),
.pxl_out(pxl_out_48), .valid_out(valid_out_48) );

//Channel 49
conv_33_s2 #(D, DATA_WIDTH) x49(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b10111111011010010001000010100100),
.kernel_01(32'b00111111011000110011001011100110),
.kernel_02(32'b10111111001110011001100110100001),
.kernel_03(32'b00111100011111110100001100101110),
.kernel_04(32'b10111110000011010110110110100001),
.kernel_05(32'b10111111100000001010010110110010),
.kernel_06(32'b10111100101000000011110100110100),
.kernel_07(32'b00111100111011000010011011110110),
.kernel_08(32'b00111111011011110110010001100000),
.pxl_out(pxl_out_49), .valid_out(valid_out_49) );

//Channel 50
conv_33_s2 #(D, DATA_WIDTH) x50(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b10111110101001100111111111011000),
.kernel_01(32'b10111110100110011101101001011111),
.kernel_02(32'b00111111000000010011011101111010),
.kernel_03(32'b10111111101010010100000001010011),
.kernel_04(32'b10111110101111011010110001010000),
.kernel_05(32'b00111111000010100010011000011000),
.kernel_06(32'b00111111000010110011001010001000),
.kernel_07(32'b10111100110001011001100111110100),
.kernel_08(32'b10111101100001111000100011001100),
.pxl_out(pxl_out_50), .valid_out(valid_out_50) );

//Channel 51
conv_33_s2 #(D, DATA_WIDTH) x51(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b00111101100010010111000100000011),
.kernel_01(32'b00111110000011001000011111101110),
.kernel_02(32'b00111101010111000000110010111110),
.kernel_03(32'b10111110111111010000010111011001),
.kernel_04(32'b00111110000100101001100001110000),
.kernel_05(32'b00111101011000101111100011001000),
.kernel_06(32'b10111011000001010001101100010101),
.kernel_07(32'b00111110100000110010110100110011),
.kernel_08(32'b10111101011110101110001010110101),
.pxl_out(pxl_out_51), .valid_out(valid_out_51) );

//Channel 52
conv_33_s2 #(D, DATA_WIDTH) x52(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b10111111010011000100101111000110),
.kernel_01(32'b00111101101111001100101001010000),
.kernel_02(32'b00111101110100101010010101100011),
.kernel_03(32'b10111101110000111001010111110110),
.kernel_04(32'b10111110001001011100100000101011),
.kernel_05(32'b00111111010010000010010100011111),
.kernel_06(32'b00111111000110001100010100001111),
.kernel_07(32'b10111100111101010000011001001000),
.kernel_08(32'b00111110000001100101000000010101),
.pxl_out(pxl_out_52), .valid_out(valid_out_52) );

//Channel 53
conv_33_s2 #(D, DATA_WIDTH) x53(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b10111110101110111100100100011001),
.kernel_01(32'b10111111001010010010010011100010),
.kernel_02(32'b00111110110011101110111000110100),
.kernel_03(32'b00111100001001000100110010011101),
.kernel_04(32'b00111111001011010000111101001101),
.kernel_05(32'b10111111010110011011010001001010),
.kernel_06(32'b10111110110001110010110101010001),
.kernel_07(32'b10111111010011000111010001011000),
.kernel_08(32'b10111111010011010010001001001001),
.pxl_out(pxl_out_53), .valid_out(valid_out_53) );

//Channel 54
conv_33_s2 #(D, DATA_WIDTH) x54(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b10111110110110100111111100111000),
.kernel_01(32'b00111110110111000100010000111101),
.kernel_02(32'b00111111000101110111101100000110),
.kernel_03(32'b00111110010000001011111101100110),
.kernel_04(32'b10111110101000101100100111011100),
.kernel_05(32'b00111110100101011000011110110110),
.kernel_06(32'b00111101110010000001111001111000),
.kernel_07(32'b00111111001101001010111001010111),
.kernel_08(32'b10111111000010001110011011101011),
.pxl_out(pxl_out_54), .valid_out(valid_out_54) );

//Channel 55
conv_33_s2 #(D, DATA_WIDTH) x55(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b00111110101000001010111011011011),
.kernel_01(32'b00111101100101110101101000010000),
.kernel_02(32'b10111110001010010010100100100010),
.kernel_03(32'b00111110001111011101101111011000),
.kernel_04(32'b10111110011100001100101001001101),
.kernel_05(32'b10111110011110001111010101100111),
.kernel_06(32'b10111110101011101001011110101110),
.kernel_07(32'b10111100010000001110011101000011),
.kernel_08(32'b00111110000101110110011010111100),
.pxl_out(pxl_out_55), .valid_out(valid_out_55) );

//Channel 56
conv_33_s2 #(D, DATA_WIDTH) x56(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b10111101111101000110001011110010),
.kernel_01(32'b00111110001010010011100000001100),
.kernel_02(32'b10111100000111101100100110000101),
.kernel_03(32'b00111110100110011100110011101110),
.kernel_04(32'b10111110100110100101000010101001),
.kernel_05(32'b00111100100110001100010000001110),
.kernel_06(32'b10111110111111000111111100101000),
.kernel_07(32'b10111110101100001110111000111011),
.kernel_08(32'b10111110110001100010100110011011),
.pxl_out(pxl_out_56), .valid_out(valid_out_56) );

//Channel 57
conv_33_s2 #(D, DATA_WIDTH) x57(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b00111111000001010101110110100110),
.kernel_01(32'b00111111001000111100111010111010),
.kernel_02(32'b00111110111101110111101110011110),
.kernel_03(32'b00111110100100100101101100111010),
.kernel_04(32'b00111111001001010010010000010101),
.kernel_05(32'b10111111000111110000101010111001),
.kernel_06(32'b10111111100001010001011110110111),
.kernel_07(32'b10111110100011010110100001101111),
.kernel_08(32'b10111101111011001101000011101101),
.pxl_out(pxl_out_57), .valid_out(valid_out_57) );

//Channel 58
conv_33_s2 #(D, DATA_WIDTH) x58(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b10111110100101010010111110111110),
.kernel_01(32'b10111100011100011010101000110111),
.kernel_02(32'b10111100111000010000100111011010),
.kernel_03(32'b00111111001111000110111101111001),
.kernel_04(32'b10111110111110100000111001000100),
.kernel_05(32'b00111110011111110001101011011001),
.kernel_06(32'b00111100110000001011010110110110),
.kernel_07(32'b00111100101100001100010001011011),
.kernel_08(32'b00111110010100111000110011110101),
.pxl_out(pxl_out_58), .valid_out(valid_out_58) );

//Channel 59
conv_33_s2 #(D, DATA_WIDTH) x59(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b00111110001010010011110111110010),
.kernel_01(32'b00111111010010110011001011000101),
.kernel_02(32'b10111110110010000110100010101111),
.kernel_03(32'b10111011101011011110001001110110),
.kernel_04(32'b10111101100111000011001100101100),
.kernel_05(32'b00111110010110010011000110010011),
.kernel_06(32'b10111111000110100000000011100111),
.kernel_07(32'b10111101000111011001001010100111),
.kernel_08(32'b10111110110101001000001000001001),
.pxl_out(pxl_out_59), .valid_out(valid_out_59) );

//Channel 60
conv_33_s2 #(D, DATA_WIDTH) x60(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b00111101101010110101011011110010),
.kernel_01(32'b00111101100000000011111101011111),
.kernel_02(32'b10111111000011111011011101100010),
.kernel_03(32'b10111101001010001011110110010100),
.kernel_04(32'b10111110111100110000110011101101),
.kernel_05(32'b00111110111111010101110100101000),
.kernel_06(32'b10111110000011000011010011101110),
.kernel_07(32'b00111111001001101000010001110010),
.kernel_08(32'b00111110001011001011101001010110),
.pxl_out(pxl_out_60), .valid_out(valid_out_60) );

//Channel 61
conv_33_s2 #(D, DATA_WIDTH) x61(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b00111111001000110001100100111001),
.kernel_01(32'b10111111000110100010100010100011),
.kernel_02(32'b10111111100100100000001100101001),
.kernel_03(32'b00111110100000011110001010011000),
.kernel_04(32'b10111100011100100100001001110100),
.kernel_05(32'b10111110101010101101111101001000),
.kernel_06(32'b00111100101000010100000101011010),
.kernel_07(32'b10111110001111101010111111101010),
.kernel_08(32'b00111110101001000111110010101101),
.pxl_out(pxl_out_61), .valid_out(valid_out_61) );

//Channel 62
conv_33_s2 #(D, DATA_WIDTH) x62(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b10111110010010010110000100001001),
.kernel_01(32'b00111110010110101100000001000100),
.kernel_02(32'b10111101010110110010100101000010),
.kernel_03(32'b00111101100100000110111110010000),
.kernel_04(32'b00111101111110100010011111100010),
.kernel_05(32'b00111110110000000101110011000110),
.kernel_06(32'b10111111000100000010111011110110),
.kernel_07(32'b10111110011110011100111101011111),
.kernel_08(32'b00111100110101011000001101100111),
.pxl_out(pxl_out_62), .valid_out(valid_out_62) );

//Channel 63
conv_33_s2 #(D, DATA_WIDTH) x63(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b10111011100100101000101110111110),
.kernel_01(32'b10111101110110110010110001000010),
.kernel_02(32'b00111110111001011000111110011010),
.kernel_03(32'b10111101100000111001101000100111),
.kernel_04(32'b00111101101001001101000010000101),
.kernel_05(32'b00111101110000010000101010001111),
.kernel_06(32'b10111101110000011001111111011101),
.kernel_07(32'b10111110101011000101001010100110),
.kernel_08(32'b00111110101010010011111110011000),
.pxl_out(pxl_out_63), .valid_out(valid_out_63) );

//Channel 64
conv_33_s2 #(D, DATA_WIDTH) x64(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b10111110001100011110011000101101),
.kernel_01(32'b00111110100100000111001101001011),
.kernel_02(32'b10111110111101010001101001111101),
.kernel_03(32'b00111110111111111101001011010000),
.kernel_04(32'b10111110110011001000011111111100),
.kernel_05(32'b00111110110100011001011010111000),
.kernel_06(32'b10111111000111110111000000001011),
.kernel_07(32'b10111111000111101111101101000011),
.kernel_08(32'b00111101110010101111001111101000),
.pxl_out(pxl_out_64), .valid_out(valid_out_64) );

//Channel 65
conv_33_s2 #(D, DATA_WIDTH) x65(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b00111110001000010110011110101110),
.kernel_01(32'b10111100011010101000011100110110),
.kernel_02(32'b00111110001000000100011110000101),
.kernel_03(32'b00111101110111100111100101000000),
.kernel_04(32'b10111111000010110110111011000110),
.kernel_05(32'b00111110111011101001110010100110),
.kernel_06(32'b10111110100001011101100111100100),
.kernel_07(32'b00111100111010110101010101001011),
.kernel_08(32'b10111101110001101111100011111001),
.pxl_out(pxl_out_65), .valid_out(valid_out_65) );

//Channel 66
conv_33_s2 #(D, DATA_WIDTH) x66(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b00111110100110001001010000000110),
.kernel_01(32'b00111110000110011100000100100111),
.kernel_02(32'b10111110000001011010111111110011),
.kernel_03(32'b10111110000010010111111101101111),
.kernel_04(32'b10111110101010000100111101100000),
.kernel_05(32'b10111110000110100111111101010110),
.kernel_06(32'b10111110001100111001000101110011),
.kernel_07(32'b00111110000110001110111000100110),
.kernel_08(32'b10111111000000010000000101100000),
.pxl_out(pxl_out_66), .valid_out(valid_out_66) );

//Channel 67
conv_33_s2 #(D, DATA_WIDTH) x67(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b00111110010011110100001011000111),
.kernel_01(32'b00111101111011010110010100111101),
.kernel_02(32'b10111101011000111110001101010010),
.kernel_03(32'b10111101011011011011010000100011),
.kernel_04(32'b10111110000001110111110110111001),
.kernel_05(32'b10111110001000100010100010011100),
.kernel_06(32'b10111111000100001100100101010110),
.kernel_07(32'b00111110110011011111010100010011),
.kernel_08(32'b10111110111000010000000111111110),
.pxl_out(pxl_out_67), .valid_out(valid_out_67) );

//Channel 68
conv_33_s2 #(D, DATA_WIDTH) x68(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b00111110011000110101001000001100),
.kernel_01(32'b00111110101001100001100010101100),
.kernel_02(32'b00111110110111011111001111011001),
.kernel_03(32'b00111110101101001100110100010011),
.kernel_04(32'b10111110100101110110011110001101),
.kernel_05(32'b10111101101100101100000001100100),
.kernel_06(32'b00111100110000111000110110000101),
.kernel_07(32'b10111101110011100011101110100010),
.kernel_08(32'b00111101101011010100100101100101),
.pxl_out(pxl_out_68), .valid_out(valid_out_68) );

//Channel 69
conv_33_s2 #(D, DATA_WIDTH) x69(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b10111111001001100100011111011100),
.kernel_01(32'b00111110111001000111101010100010),
.kernel_02(32'b10111110001011110010011110011001),
.kernel_03(32'b00111110000010100101101011110011),
.kernel_04(32'b10111101100011100000100011110110),
.kernel_05(32'b00111110110110100110111010011001),
.kernel_06(32'b00111101100001010101001001111000),
.kernel_07(32'b00111110111100000101011011011001),
.kernel_08(32'b10111101100110001100010010111111),
.pxl_out(pxl_out_69), .valid_out(valid_out_69) );

//Channel 70
conv_33_s2 #(D, DATA_WIDTH) x70(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b10111110111100101001011011010011),
.kernel_01(32'b00111100101001000110001001010010),
.kernel_02(32'b00111110001011001001101010010010),
.kernel_03(32'b10111110110010101010110011010110),
.kernel_04(32'b10111110101110100000001011110001),
.kernel_05(32'b10111110100000100110011011101100),
.kernel_06(32'b10111101101110000110100001110100),
.kernel_07(32'b10111100100000110000000111111001),
.kernel_08(32'b00111010111000011111011101111110),
.pxl_out(pxl_out_70), .valid_out(valid_out_70) );

//Channel 71
conv_33_s2 #(D, DATA_WIDTH) x71(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b00111101110000100100101100110101),
.kernel_01(32'b10111110011110001011000101110000),
.kernel_02(32'b10111111000001000111100100011111),
.kernel_03(32'b10111101101110001001010101000111),
.kernel_04(32'b10111110110111110010011100100001),
.kernel_05(32'b00111110000001110101111010100010),
.kernel_06(32'b00111110110001111000100011100000),
.kernel_07(32'b00111111000000001100001101011000),
.kernel_08(32'b00111110110011001011101010011101),
.pxl_out(pxl_out_71), .valid_out(valid_out_71) );

//Channel 72
conv_33_s2 #(D, DATA_WIDTH) x72(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b00111110001101001001100111000001),
.kernel_01(32'b10111101010111011001111101000000),
.kernel_02(32'b00111101101110101110010111100001),
.kernel_03(32'b10111101001011100101001010001111),
.kernel_04(32'b00111101010001110001100010110001),
.kernel_05(32'b10111110101011011101110101010100),
.kernel_06(32'b00111110010100100011001000101011),
.kernel_07(32'b00111110000010110101111011010001),
.kernel_08(32'b00111110010011100110010110110011),
.pxl_out(pxl_out_72), .valid_out(valid_out_72) );

//Channel 73
conv_33_s2 #(D, DATA_WIDTH) x73(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b00111100110011110011010100111000),
.kernel_01(32'b00111101111110011111100010110011),
.kernel_02(32'b10111110011010110110110000001000),
.kernel_03(32'b10111110101101100101110110010010),
.kernel_04(32'b10111101100110100000001010001010),
.kernel_05(32'b10111110011110101001100001001111),
.kernel_06(32'b00111101100111100000110010011111),
.kernel_07(32'b10111101010001000000101110001000),
.kernel_08(32'b00111110011111101011101111110001),
.pxl_out(pxl_out_73), .valid_out(valid_out_73) );

//Channel 74
conv_33_s2 #(D, DATA_WIDTH) x74(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b10111110010110011111100001101100),
.kernel_01(32'b00111101000110010000110001001100),
.kernel_02(32'b10111101010110011111000010000000),
.kernel_03(32'b10111101010000000110011111111000),
.kernel_04(32'b10111100101111001010100111101010),
.kernel_05(32'b00111110010010000001110010111010),
.kernel_06(32'b10111110001010000011111011001011),
.kernel_07(32'b10111110100000001100110110011111),
.kernel_08(32'b10111110101111100010110100001001),
.pxl_out(pxl_out_74), .valid_out(valid_out_74) );

//Channel 75
conv_33_s2 #(D, DATA_WIDTH) x75(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b10111110110110110000110101100000),
.kernel_01(32'b10111110100010000110001011001001),
.kernel_02(32'b00111110100000110001011110111001),
.kernel_03(32'b00111110110010010111111001001111),
.kernel_04(32'b00111110001010100010011011001010),
.kernel_05(32'b00111110000010000010111010011100),
.kernel_06(32'b00111101011110110000101111101010),
.kernel_07(32'b10111100111110100001110001010010),
.kernel_08(32'b00111110100011001100111111100010),
.pxl_out(pxl_out_75), .valid_out(valid_out_75) );

//Channel 76
conv_33_s2 #(D, DATA_WIDTH) x76(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b00111110001010100110010110100010),
.kernel_01(32'b10111101000001100111011000010011),
.kernel_02(32'b00111111011101010000001111010001),
.kernel_03(32'b10111110001000011101001000011101),
.kernel_04(32'b00111101010111000100111110010000),
.kernel_05(32'b10111110010000110011001101100001),
.kernel_06(32'b00111111001110100010010111101000),
.kernel_07(32'b00111100011011010101110010001111),
.kernel_08(32'b10111110100000101110111001110010),
.pxl_out(pxl_out_76), .valid_out(valid_out_76) );

//Channel 77
conv_33_s2 #(D, DATA_WIDTH) x77(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b00111101000010011100001110011101),
.kernel_01(32'b10111111011101011010000111100011),
.kernel_02(32'b10111110101110001010101100100101),
.kernel_03(32'b10111110101000010010110010110101),
.kernel_04(32'b00111110011000000000100110100000),
.kernel_05(32'b00111111000101100000101001001111),
.kernel_06(32'b00111110100011111101000101111111),
.kernel_07(32'b10111101110100011111010100110110),
.kernel_08(32'b00111101101001110100100000100110),
.pxl_out(pxl_out_77), .valid_out(valid_out_77) );

//Channel 78
conv_33_s2 #(D, DATA_WIDTH) x78(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b10111101010000011111010000000000),
.kernel_01(32'b10111110011101111111010000010100),
.kernel_02(32'b10111101100111100000101111101001),
.kernel_03(32'b10111111010111110000110110110101),
.kernel_04(32'b00111111001000110100000110011101),
.kernel_05(32'b10111110100110111000111001100011),
.kernel_06(32'b00111110110011100111000100001011),
.kernel_07(32'b10111111010010110101111101011110),
.kernel_08(32'b10111110101000000000110011011000),
.pxl_out(pxl_out_78), .valid_out(valid_out_78) );

//Channel 79
conv_33_s2 #(D, DATA_WIDTH) x79(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b00111110111011010101010110011111),
.kernel_01(32'b10111110111111011011101000010100),
.kernel_02(32'b10111101010010000111101111000110),
.kernel_03(32'b00111100001100100110111101101000),
.kernel_04(32'b10111101111000000001111111110110),
.kernel_05(32'b00111100111111101011011111010100),
.kernel_06(32'b10111011010011101000100100100101),
.kernel_07(32'b00111111100000111101010010000101),
.kernel_08(32'b10111101100101010000100101010111),
.pxl_out(pxl_out_79), .valid_out(valid_out_79) );

//Channel 80
conv_33_s2 #(D, DATA_WIDTH) x80(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b00111110011000001000101111000110),
.kernel_01(32'b10111110000110000011011010011111),
.kernel_02(32'b00111111011101111000111110000011),
.kernel_03(32'b00111110000111001011111101000110),
.kernel_04(32'b00111111010001011000010111000000),
.kernel_05(32'b00111101001011110001101100101011),
.kernel_06(32'b10111111100111111101111101001011),
.kernel_07(32'b10111110000010000100000111011111),
.kernel_08(32'b00111110100100011100010101011110),
.pxl_out(pxl_out_80), .valid_out(valid_out_80) );

//Channel 81
conv_33_s2 #(D, DATA_WIDTH) x81(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b10111111000111111100001110110000),
.kernel_01(32'b00111110111100000000100110001101),
.kernel_02(32'b10111110101111010110011010111101),
.kernel_03(32'b10111101010010100010000101001000),
.kernel_04(32'b00111101001100100000110101000011),
.kernel_05(32'b10111101100111011100000010011111),
.kernel_06(32'b00111100110000000101101000011010),
.kernel_07(32'b10111110000001111100100101111010),
.kernel_08(32'b10111111011010011110101111001001),
.pxl_out(pxl_out_81), .valid_out(valid_out_81) );

//Channel 82
conv_33_s2 #(D, DATA_WIDTH) x82(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b10111110001000101011000111000010),
.kernel_01(32'b10111110001111101111011000110011),
.kernel_02(32'b00111110100010000101101100111011),
.kernel_03(32'b10111111001101010001010110100100),
.kernel_04(32'b10111110010000100010110101110000),
.kernel_05(32'b00111110111000111111100001111010),
.kernel_06(32'b00111110101001101011100001100111),
.kernel_07(32'b10111100101001110011101010001101),
.kernel_08(32'b00111101000110011010111111110000),
.pxl_out(pxl_out_82), .valid_out(valid_out_82) );

//Channel 83
conv_33_s2 #(D, DATA_WIDTH) x83(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b10111101010111111011101111000000),
.kernel_01(32'b10111101000011011001100100011101),
.kernel_02(32'b00111100110001100100010000101100),
.kernel_03(32'b00111111001010110010010001010010),
.kernel_04(32'b00111101001111101000011100111111),
.kernel_05(32'b00111110111100111011111101011001),
.kernel_06(32'b10111101101111001000010010110100),
.kernel_07(32'b00111110111100110000011101010111),
.kernel_08(32'b10111101101101010011011011011111),
.pxl_out(pxl_out_83), .valid_out(valid_out_83) );

//Channel 84
conv_33_s2 #(D, DATA_WIDTH) x84(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b10111111000011001100010100001111),
.kernel_01(32'b00111101011000111100011100000000),
.kernel_02(32'b10111111001000100100101011100000),
.kernel_03(32'b10111101110010111100010100001111),
.kernel_04(32'b10111110000001001011101101101100),
.kernel_05(32'b00111110110001101111111110101000),
.kernel_06(32'b00111110100100001001101101001110),
.kernel_07(32'b00111101111111110000110100000011),
.kernel_08(32'b00111101100111000011111110010001),
.pxl_out(pxl_out_84), .valid_out(valid_out_84) );

//Channel 85
conv_33_s2 #(D, DATA_WIDTH) x85(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b10111101110110001101010101000111),
.kernel_01(32'b10111110000001000001101110101010),
.kernel_02(32'b00111110100100100100001111111100),
.kernel_03(32'b10111101010001111111111000000101),
.kernel_04(32'b10111111000001110111100001100111),
.kernel_05(32'b10111111000000111011001111001011),
.kernel_06(32'b10111110010000101010101000010000),
.kernel_07(32'b10111110111001110001110011010010),
.kernel_08(32'b10111110101001111101011010110010),
.pxl_out(pxl_out_85), .valid_out(valid_out_85) );

//Channel 86
conv_33_s2 #(D, DATA_WIDTH) x86(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b10111110001101101110110101101101),
.kernel_01(32'b00111110100010111100001011101011),
.kernel_02(32'b00111110100001001011001011000100),
.kernel_03(32'b00111110001111011110011101101111),
.kernel_04(32'b10111101101111100100110000011100),
.kernel_05(32'b00111110011010011111001111001111),
.kernel_06(32'b00111101100100001000011011001101),
.kernel_07(32'b00111111000101100101010001111100),
.kernel_08(32'b00111110110111011011100000110101),
.pxl_out(pxl_out_86), .valid_out(valid_out_86) );

//Channel 87
conv_33_s2 #(D, DATA_WIDTH) x87(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b00111101100000011111111111111001),
.kernel_01(32'b00111101011011110000011100101010),
.kernel_02(32'b10111101100011001111000110011011),
.kernel_03(32'b00111110100001101001011001110000),
.kernel_04(32'b10111110001010000110010010110010),
.kernel_05(32'b10111110000101001110011001000101),
.kernel_06(32'b00111101011001010001100100011100),
.kernel_07(32'b10111111000001010000101001110100),
.kernel_08(32'b10111110100100001111011111001111),
.pxl_out(pxl_out_87), .valid_out(valid_out_87) );

//Channel 88
conv_33_s2 #(D, DATA_WIDTH) x88(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b10111101101100000110110010010101),
.kernel_01(32'b00111110000100100110110111011010),
.kernel_02(32'b10111101101100110101101100011011),
.kernel_03(32'b00111101000000100111000011001000),
.kernel_04(32'b10111101001101001100110110100010),
.kernel_05(32'b10111011100011000110111001000100),
.kernel_06(32'b10111011111111011111011110010110),
.kernel_07(32'b10111110100001001111001111011110),
.kernel_08(32'b00111110001011110011000111111000),
.pxl_out(pxl_out_88), .valid_out(valid_out_88) );

//Channel 89
conv_33_s2 #(D, DATA_WIDTH) x89(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b10111111000010110000011010100011),
.kernel_01(32'b00111110110001011011000101010011),
.kernel_02(32'b00111110101010001100111011000001),
.kernel_03(32'b00111110011000010101011100111100),
.kernel_04(32'b00111110101100010011001000011000),
.kernel_05(32'b10111110101111111111110010010100),
.kernel_06(32'b10111111001111110101110010101110),
.kernel_07(32'b10111110001011000000110110100011),
.kernel_08(32'b10111110000001111001100001010101),
.pxl_out(pxl_out_89), .valid_out(valid_out_89) );

//Channel 90
conv_33_s2 #(D, DATA_WIDTH) x90(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b00111100111101010001100100100101),
.kernel_01(32'b10111100101000111100010010111011),
.kernel_02(32'b10111101011111110101011011000100),
.kernel_03(32'b00111111001011110111101100100001),
.kernel_04(32'b00111110111001111110010100101100),
.kernel_05(32'b00111101011001110010011100110101),
.kernel_06(32'b00111110000011010111010011010110),
.kernel_07(32'b10111011111011100010111000000101),
.kernel_08(32'b00111110111110100100001000001110),
.pxl_out(pxl_out_90), .valid_out(valid_out_90) );

//Channel 91
conv_33_s2 #(D, DATA_WIDTH) x91(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b00111110001100000011101101011101),
.kernel_01(32'b00111110111111100100111100010100),
.kernel_02(32'b00111101001000110101000011111110),
.kernel_03(32'b10111111001100011111001101111010),
.kernel_04(32'b00111101001001111011110111101110),
.kernel_05(32'b00111110000111011001101110000111),
.kernel_06(32'b10111110101110101000001101101011),
.kernel_07(32'b10111110000001101100001010001011),
.kernel_08(32'b10111101111110001001101110000100),
.pxl_out(pxl_out_91), .valid_out(valid_out_91) );

//Channel 92
conv_33_s2 #(D, DATA_WIDTH) x92(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b00111100001000111111011001001111),
.kernel_01(32'b00111101000001111100001001011010),
.kernel_02(32'b00111011110111010000100010110111),
.kernel_03(32'b10111100001101101000011010111100),
.kernel_04(32'b00111110100110000000001011111111),
.kernel_05(32'b10111111000000010110011010011011),
.kernel_06(32'b10111101101011101000111000111110),
.kernel_07(32'b00111110110101000111001111101111),
.kernel_08(32'b00111101101000100100100100100110),
.pxl_out(pxl_out_92), .valid_out(valid_out_92) );

//Channel 93
conv_33_s2 #(D, DATA_WIDTH) x93(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b00111110101100011001011111000100),
.kernel_01(32'b10111110101100100100001100101110),
.kernel_02(32'b10111111010100100010000010011100),
.kernel_03(32'b00111110001000100001100001110001),
.kernel_04(32'b10111100001100001000000001001100),
.kernel_05(32'b10111100011001111010011111111110),
.kernel_06(32'b10111101010101010011100001101111),
.kernel_07(32'b10111110001011011101111000101001),
.kernel_08(32'b00111110101010011111001101010101),
.pxl_out(pxl_out_93), .valid_out(valid_out_93) );

//Channel 94
conv_33_s2 #(D, DATA_WIDTH) x94(.clk(clk), .reset(reset), .valid_in(valid_in_1), .pxl_in(pxl_in_1),
.kernel_00(32'b00111110011101011101110011000001),
.kernel_01(32'b00111101001011110000011010110011),
.kernel_02(32'b00111110001110100010000110111001),
.kernel_03(32'b00111010101101111001011101011000),
.kernel_04(32'b00111110011000011101000101001010),
.kernel_05(32'b00111110001000000011111010110010),
.kernel_06(32'b10111110101110110111111011001001),
.kernel_07(32'b00111101101011001101001101111011),
.kernel_08(32'b10111110101111011111101001010110),
.pxl_out(pxl_out_94), .valid_out(valid_out_94) );

//Channel 95
conv_33_s2 #(D, DATA_WIDTH) x95(.clk(clk), .reset(reset), .valid_in(valid_in_2), .pxl_in(pxl_in_2),
.kernel_00(32'b00111101101001111000010010101110),
.kernel_01(32'b10111101011111100111001000001101),
.kernel_02(32'b00111110010110111011011111011000),
.kernel_03(32'b10111101110010011010011110010010),
.kernel_04(32'b00111101111010001000110110011001),
.kernel_05(32'b00111101000000001001101000010110),
.kernel_06(32'b00111100000100001101100101011110),
.kernel_07(32'b10111101000000100010001001011101),
.kernel_08(32'b00111110010001101111100010101001),
.pxl_out(pxl_out_95), .valid_out(valid_out_95) );

//Channel 96
conv_33_s2 #(D, DATA_WIDTH) x96(.clk(clk), .reset(reset), .valid_in(valid_in_3), .pxl_in(pxl_in_3),
.kernel_00(32'b00111110010000010100011010000101),
.kernel_01(32'b10111110011011100101101000101101),
.kernel_02(32'b10111110100110100101000010001001),
.kernel_03(32'b00111110101110010100100001010110),
.kernel_04(32'b10111110010001000001001110010000),
.kernel_05(32'b00111110010011101000010110101001),
.kernel_06(32'b10111110101011000000011100010011),
.kernel_07(32'b10111110111000010010001010100100),
.kernel_08(32'b00111100111001000000100100010000),
.pxl_out(pxl_out_96), .valid_out(valid_out_96) );


endmodule