// Convolution Kernel 3x3, Stride = 1, Padding = 0, Channel = 32.
//Input = 149x149x32, Output = 147x147x32.

module CONV_3x3_Stride1_32
#(parameter D = 220,
  parameter DATA_WIDTH = 32)
(
     //input
    	input clk,
     	input reset,
     	input valid_in_1,valid_in_2,valid_in_3,valid_in_4,valid_in_5,valid_in_6,valid_in_7,valid_in_8,valid_in_9,
            valid_in_10,valid_in_11,valid_in_12,valid_in_13,valid_in_14,valid_in_15,valid_in_16,valid_in_17,valid_in_18,
            valid_in_19,valid_in_20,valid_in_21,valid_in_22,valid_in_23,valid_in_24,valid_in_25,valid_in_26,valid_in_27,
            valid_in_28,valid_in_29,valid_in_30,valid_in_31,valid_in_32,
            
      input [DATA_WIDTH-1:0] pxl_in_1,pxl_in_2,pxl_in_3,pxl_in_4,pxl_in_5,pxl_in_6,pxl_in_7,pxl_in_8,pxl_in_9,
                             pxl_in_10,pxl_in_11,pxl_in_12,pxl_in_13,pxl_in_14,pxl_in_15,pxl_in_16,pxl_in_17,pxl_in_18,
                             pxl_in_19,pxl_in_20,pxl_in_21,pxl_in_22,pxl_in_23,pxl_in_24,pxl_in_25,pxl_in_26,pxl_in_27,
                             pxl_in_28,pxl_in_29,pxl_in_30,pxl_in_31,pxl_in_32,
    
     output [DATA_WIDTH-1:0] pxl_out_1 , pxl_out_2 , pxl_out_3 , pxl_out_4 , pxl_out_5 , pxl_out_6 , pxl_out_7 , pxl_out_8 , pxl_out_9 , pxl_out_10,
                        pxl_out_11, pxl_out_12, pxl_out_13, pxl_out_14, pxl_out_15, pxl_out_16, pxl_out_17, pxl_out_18, pxl_out_19, pxl_out_20,
	                      pxl_out_21, pxl_out_22, pxl_out_23, pxl_out_24, pxl_out_25, pxl_out_26, pxl_out_27, pxl_out_28, pxl_out_29, pxl_out_30,
                        pxl_out_31, pxl_out_32,
	                                 
	               output valid_out_1 , valid_out_2 , valid_out_3 , valid_out_4 , valid_out_5 , valid_out_6 , valid_out_7 , valid_out_8 , valid_out_9 , valid_out_10,
                        valid_out_11, valid_out_12, valid_out_13, valid_out_14, valid_out_15, valid_out_16, valid_out_17, valid_out_18, valid_out_19, valid_out_20,
	                      valid_out_21, valid_out_22, valid_out_23, valid_out_24, valid_out_25, valid_out_26, valid_out_27, valid_out_28, valid_out_29, valid_out_30,
                        valid_out_31, valid_out_32
                        
);
wire [DATA_WIDTH-1:0] tmp_pxl_out_1, tmp_pxl_out_2, tmp_pxl_out_3, tmp_pxl_out_4, tmp_pxl_out_5, tmp_pxl_out_6, tmp_pxl_out_7, tmp_pxl_out_8, tmp_pxl_out_9, 
tmp_pxl_out_10, tmp_pxl_out_11, tmp_pxl_out_12, tmp_pxl_out_13, tmp_pxl_out_14, tmp_pxl_out_15, tmp_pxl_out_16, tmp_pxl_out_17, tmp_pxl_out_18, 
tmp_pxl_out_19, tmp_pxl_out_20, tmp_pxl_out_21, tmp_pxl_out_22, tmp_pxl_out_23, tmp_pxl_out_24, tmp_pxl_out_25, tmp_pxl_out_26, tmp_pxl_out_27, 
tmp_pxl_out_28, tmp_pxl_out_29, tmp_pxl_out_30, tmp_pxl_out_31, tmp_pxl_out_32, tmp_pxl_out_33, tmp_pxl_out_34, tmp_pxl_out_35, tmp_pxl_out_36, 
tmp_pxl_out_37, tmp_pxl_out_38, tmp_pxl_out_39, tmp_pxl_out_40, tmp_pxl_out_41, tmp_pxl_out_42, tmp_pxl_out_43, tmp_pxl_out_44, tmp_pxl_out_45, 
tmp_pxl_out_46, tmp_pxl_out_47, tmp_pxl_out_48, tmp_pxl_out_49, tmp_pxl_out_50, tmp_pxl_out_51, tmp_pxl_out_52, tmp_pxl_out_53, tmp_pxl_out_54, 
tmp_pxl_out_55, tmp_pxl_out_56, tmp_pxl_out_57, tmp_pxl_out_58, tmp_pxl_out_59, tmp_pxl_out_60, tmp_pxl_out_61, tmp_pxl_out_62, tmp_pxl_out_63, 
tmp_pxl_out_64, tmp_pxl_out_65, tmp_pxl_out_66, tmp_pxl_out_67, tmp_pxl_out_68, tmp_pxl_out_69, tmp_pxl_out_70, tmp_pxl_out_71, tmp_pxl_out_72, 
tmp_pxl_out_73, tmp_pxl_out_74, tmp_pxl_out_75, tmp_pxl_out_76, tmp_pxl_out_77, tmp_pxl_out_78, tmp_pxl_out_79, tmp_pxl_out_80, tmp_pxl_out_81, 
tmp_pxl_out_82, tmp_pxl_out_83, tmp_pxl_out_84, tmp_pxl_out_85, tmp_pxl_out_86, tmp_pxl_out_87, tmp_pxl_out_88, tmp_pxl_out_89, tmp_pxl_out_90, 
tmp_pxl_out_91, tmp_pxl_out_92, tmp_pxl_out_93, tmp_pxl_out_94, tmp_pxl_out_95, tmp_pxl_out_96, tmp_pxl_out_97, tmp_pxl_out_98, tmp_pxl_out_99, 
tmp_pxl_out_100, tmp_pxl_out_101, tmp_pxl_out_102, tmp_pxl_out_103, tmp_pxl_out_104, tmp_pxl_out_105, tmp_pxl_out_106, tmp_pxl_out_107, tmp_pxl_out_108, 
tmp_pxl_out_109, tmp_pxl_out_110, tmp_pxl_out_111, tmp_pxl_out_112, tmp_pxl_out_113, tmp_pxl_out_114, tmp_pxl_out_115, tmp_pxl_out_116, tmp_pxl_out_117, 
tmp_pxl_out_118, tmp_pxl_out_119, tmp_pxl_out_120, tmp_pxl_out_121, tmp_pxl_out_122, tmp_pxl_out_123, tmp_pxl_out_124, tmp_pxl_out_125, tmp_pxl_out_126, 
tmp_pxl_out_127, tmp_pxl_out_128, tmp_pxl_out_129, tmp_pxl_out_130, tmp_pxl_out_131, tmp_pxl_out_132, tmp_pxl_out_133, tmp_pxl_out_134, tmp_pxl_out_135, 
tmp_pxl_out_136, tmp_pxl_out_137, tmp_pxl_out_138, tmp_pxl_out_139, tmp_pxl_out_140, tmp_pxl_out_141, tmp_pxl_out_142, tmp_pxl_out_143, tmp_pxl_out_144, 
tmp_pxl_out_145, tmp_pxl_out_146, tmp_pxl_out_147, tmp_pxl_out_148, tmp_pxl_out_149, tmp_pxl_out_150, tmp_pxl_out_151, tmp_pxl_out_152, tmp_pxl_out_153, 
tmp_pxl_out_154, tmp_pxl_out_155, tmp_pxl_out_156, tmp_pxl_out_157, tmp_pxl_out_158, tmp_pxl_out_159, tmp_pxl_out_160, tmp_pxl_out_161, tmp_pxl_out_162, 
tmp_pxl_out_163, tmp_pxl_out_164, tmp_pxl_out_165, tmp_pxl_out_166, tmp_pxl_out_167, tmp_pxl_out_168, tmp_pxl_out_169, tmp_pxl_out_170, tmp_pxl_out_171, 
tmp_pxl_out_172, tmp_pxl_out_173, tmp_pxl_out_174, tmp_pxl_out_175, tmp_pxl_out_176, tmp_pxl_out_177, tmp_pxl_out_178, tmp_pxl_out_179, tmp_pxl_out_180, 
tmp_pxl_out_181, tmp_pxl_out_182, tmp_pxl_out_183, tmp_pxl_out_184, tmp_pxl_out_185, tmp_pxl_out_186, tmp_pxl_out_187, tmp_pxl_out_188, tmp_pxl_out_189, 
tmp_pxl_out_190, tmp_pxl_out_191, tmp_pxl_out_192, tmp_pxl_out_193, tmp_pxl_out_194, tmp_pxl_out_195, tmp_pxl_out_196, tmp_pxl_out_197, tmp_pxl_out_198, 
tmp_pxl_out_199, tmp_pxl_out_200, tmp_pxl_out_201, tmp_pxl_out_202, tmp_pxl_out_203, tmp_pxl_out_204, tmp_pxl_out_205, tmp_pxl_out_206, tmp_pxl_out_207, 
tmp_pxl_out_208, tmp_pxl_out_209, tmp_pxl_out_210, tmp_pxl_out_211, tmp_pxl_out_212, tmp_pxl_out_213, tmp_pxl_out_214, tmp_pxl_out_215, tmp_pxl_out_216, 
tmp_pxl_out_217, tmp_pxl_out_218, tmp_pxl_out_219, tmp_pxl_out_220, tmp_pxl_out_221, tmp_pxl_out_222, tmp_pxl_out_223, tmp_pxl_out_224, tmp_pxl_out_225, 
tmp_pxl_out_226, tmp_pxl_out_227, tmp_pxl_out_228, tmp_pxl_out_229, tmp_pxl_out_230, tmp_pxl_out_231, tmp_pxl_out_232, tmp_pxl_out_233, tmp_pxl_out_234, 
tmp_pxl_out_235, tmp_pxl_out_236, tmp_pxl_out_237, tmp_pxl_out_238, tmp_pxl_out_239, tmp_pxl_out_240, tmp_pxl_out_241, tmp_pxl_out_242, tmp_pxl_out_243, 
tmp_pxl_out_244, tmp_pxl_out_245, tmp_pxl_out_246, tmp_pxl_out_247, tmp_pxl_out_248, tmp_pxl_out_249, tmp_pxl_out_250, tmp_pxl_out_251, tmp_pxl_out_252, 
tmp_pxl_out_253, tmp_pxl_out_254, tmp_pxl_out_255, tmp_pxl_out_256, tmp_pxl_out_257, tmp_pxl_out_258, tmp_pxl_out_259, tmp_pxl_out_260, tmp_pxl_out_261, 
tmp_pxl_out_262, tmp_pxl_out_263, tmp_pxl_out_264, tmp_pxl_out_265, tmp_pxl_out_266, tmp_pxl_out_267, tmp_pxl_out_268, tmp_pxl_out_269, tmp_pxl_out_270, 
tmp_pxl_out_271, tmp_pxl_out_272, tmp_pxl_out_273, tmp_pxl_out_274, tmp_pxl_out_275, tmp_pxl_out_276, tmp_pxl_out_277, tmp_pxl_out_278, tmp_pxl_out_279, 
tmp_pxl_out_280, tmp_pxl_out_281, tmp_pxl_out_282, tmp_pxl_out_283, tmp_pxl_out_284, tmp_pxl_out_285, tmp_pxl_out_286, tmp_pxl_out_287, tmp_pxl_out_288, 
tmp_pxl_out_289, tmp_pxl_out_290, tmp_pxl_out_291, tmp_pxl_out_292, tmp_pxl_out_293, tmp_pxl_out_294, tmp_pxl_out_295, tmp_pxl_out_296, tmp_pxl_out_297, 
tmp_pxl_out_298, tmp_pxl_out_299, tmp_pxl_out_300, tmp_pxl_out_301, tmp_pxl_out_302, tmp_pxl_out_303, tmp_pxl_out_304, tmp_pxl_out_305, tmp_pxl_out_306, 
tmp_pxl_out_307, tmp_pxl_out_308, tmp_pxl_out_309, tmp_pxl_out_310, tmp_pxl_out_311, tmp_pxl_out_312, tmp_pxl_out_313, tmp_pxl_out_314, tmp_pxl_out_315, 
tmp_pxl_out_316, tmp_pxl_out_317, tmp_pxl_out_318, tmp_pxl_out_319, tmp_pxl_out_320, tmp_pxl_out_321, tmp_pxl_out_322, tmp_pxl_out_323, tmp_pxl_out_324, 
tmp_pxl_out_325, tmp_pxl_out_326, tmp_pxl_out_327, tmp_pxl_out_328, tmp_pxl_out_329, tmp_pxl_out_330, tmp_pxl_out_331, tmp_pxl_out_332, tmp_pxl_out_333, 
tmp_pxl_out_334, tmp_pxl_out_335, tmp_pxl_out_336, tmp_pxl_out_337, tmp_pxl_out_338, tmp_pxl_out_339, tmp_pxl_out_340, tmp_pxl_out_341, tmp_pxl_out_342, 
tmp_pxl_out_343, tmp_pxl_out_344, tmp_pxl_out_345, tmp_pxl_out_346, tmp_pxl_out_347, tmp_pxl_out_348, tmp_pxl_out_349, tmp_pxl_out_350, tmp_pxl_out_351, 
tmp_pxl_out_352, tmp_pxl_out_353, tmp_pxl_out_354, tmp_pxl_out_355, tmp_pxl_out_356, tmp_pxl_out_357, tmp_pxl_out_358, tmp_pxl_out_359, tmp_pxl_out_360, 
tmp_pxl_out_361, tmp_pxl_out_362, tmp_pxl_out_363, tmp_pxl_out_364, tmp_pxl_out_365, tmp_pxl_out_366, tmp_pxl_out_367, tmp_pxl_out_368, tmp_pxl_out_369, 
tmp_pxl_out_370, tmp_pxl_out_371, tmp_pxl_out_372, tmp_pxl_out_373, tmp_pxl_out_374, tmp_pxl_out_375, tmp_pxl_out_376, tmp_pxl_out_377, tmp_pxl_out_378, 
tmp_pxl_out_379, tmp_pxl_out_380, tmp_pxl_out_381, tmp_pxl_out_382, tmp_pxl_out_383, tmp_pxl_out_384, tmp_pxl_out_385, tmp_pxl_out_386, tmp_pxl_out_387, 
tmp_pxl_out_388, tmp_pxl_out_389, tmp_pxl_out_390, tmp_pxl_out_391, tmp_pxl_out_392, tmp_pxl_out_393, tmp_pxl_out_394, tmp_pxl_out_395, tmp_pxl_out_396, 
tmp_pxl_out_397, tmp_pxl_out_398, tmp_pxl_out_399, tmp_pxl_out_400, tmp_pxl_out_401, tmp_pxl_out_402, tmp_pxl_out_403, tmp_pxl_out_404, tmp_pxl_out_405, 
tmp_pxl_out_406, tmp_pxl_out_407, tmp_pxl_out_408, tmp_pxl_out_409, tmp_pxl_out_410, tmp_pxl_out_411, tmp_pxl_out_412, tmp_pxl_out_413, tmp_pxl_out_414, 
tmp_pxl_out_415, tmp_pxl_out_416, tmp_pxl_out_417, tmp_pxl_out_418, tmp_pxl_out_419, tmp_pxl_out_420, tmp_pxl_out_421, tmp_pxl_out_422, tmp_pxl_out_423, 
tmp_pxl_out_424, tmp_pxl_out_425, tmp_pxl_out_426, tmp_pxl_out_427, tmp_pxl_out_428, tmp_pxl_out_429, tmp_pxl_out_430, tmp_pxl_out_431, tmp_pxl_out_432, 
tmp_pxl_out_433, tmp_pxl_out_434, tmp_pxl_out_435, tmp_pxl_out_436, tmp_pxl_out_437, tmp_pxl_out_438, tmp_pxl_out_439, tmp_pxl_out_440, tmp_pxl_out_441, 
tmp_pxl_out_442, tmp_pxl_out_443, tmp_pxl_out_444, tmp_pxl_out_445, tmp_pxl_out_446, tmp_pxl_out_447, tmp_pxl_out_448, tmp_pxl_out_449, tmp_pxl_out_450, 
tmp_pxl_out_451, tmp_pxl_out_452, tmp_pxl_out_453, tmp_pxl_out_454, tmp_pxl_out_455, tmp_pxl_out_456, tmp_pxl_out_457, tmp_pxl_out_458, tmp_pxl_out_459, 
tmp_pxl_out_460, tmp_pxl_out_461, tmp_pxl_out_462, tmp_pxl_out_463, tmp_pxl_out_464, tmp_pxl_out_465, tmp_pxl_out_466, tmp_pxl_out_467, tmp_pxl_out_468, 
tmp_pxl_out_469, tmp_pxl_out_470, tmp_pxl_out_471, tmp_pxl_out_472, tmp_pxl_out_473, tmp_pxl_out_474, tmp_pxl_out_475, tmp_pxl_out_476, tmp_pxl_out_477, 
tmp_pxl_out_478, tmp_pxl_out_479, tmp_pxl_out_480, tmp_pxl_out_481, tmp_pxl_out_482, tmp_pxl_out_483, tmp_pxl_out_484, tmp_pxl_out_485, tmp_pxl_out_486, 
tmp_pxl_out_487, tmp_pxl_out_488, tmp_pxl_out_489, tmp_pxl_out_490, tmp_pxl_out_491, tmp_pxl_out_492, tmp_pxl_out_493, tmp_pxl_out_494, tmp_pxl_out_495, 
tmp_pxl_out_496, tmp_pxl_out_497, tmp_pxl_out_498, tmp_pxl_out_499, tmp_pxl_out_500, tmp_pxl_out_501, tmp_pxl_out_502, tmp_pxl_out_503, tmp_pxl_out_504, 
tmp_pxl_out_505, tmp_pxl_out_506, tmp_pxl_out_507, tmp_pxl_out_508, tmp_pxl_out_509, tmp_pxl_out_510, tmp_pxl_out_511, tmp_pxl_out_512, tmp_pxl_out_513, 
tmp_pxl_out_514, tmp_pxl_out_515, tmp_pxl_out_516, tmp_pxl_out_517, tmp_pxl_out_518, tmp_pxl_out_519, tmp_pxl_out_520, tmp_pxl_out_521, tmp_pxl_out_522, 
tmp_pxl_out_523, tmp_pxl_out_524, tmp_pxl_out_525, tmp_pxl_out_526, tmp_pxl_out_527, tmp_pxl_out_528, tmp_pxl_out_529, tmp_pxl_out_530, tmp_pxl_out_531, 
tmp_pxl_out_532, tmp_pxl_out_533, tmp_pxl_out_534, tmp_pxl_out_535, tmp_pxl_out_536, tmp_pxl_out_537, tmp_pxl_out_538, tmp_pxl_out_539, tmp_pxl_out_540, 
tmp_pxl_out_541, tmp_pxl_out_542, tmp_pxl_out_543, tmp_pxl_out_544, tmp_pxl_out_545, tmp_pxl_out_546, tmp_pxl_out_547, tmp_pxl_out_548, tmp_pxl_out_549, 
tmp_pxl_out_550, tmp_pxl_out_551, tmp_pxl_out_552, tmp_pxl_out_553, tmp_pxl_out_554, tmp_pxl_out_555, tmp_pxl_out_556, tmp_pxl_out_557, tmp_pxl_out_558, 
tmp_pxl_out_559, tmp_pxl_out_560, tmp_pxl_out_561, tmp_pxl_out_562, tmp_pxl_out_563, tmp_pxl_out_564, tmp_pxl_out_565, tmp_pxl_out_566, tmp_pxl_out_567, 
tmp_pxl_out_568, tmp_pxl_out_569, tmp_pxl_out_570, tmp_pxl_out_571, tmp_pxl_out_572, tmp_pxl_out_573, tmp_pxl_out_574, tmp_pxl_out_575, tmp_pxl_out_576, 
tmp_pxl_out_577, tmp_pxl_out_578, tmp_pxl_out_579, tmp_pxl_out_580, tmp_pxl_out_581, tmp_pxl_out_582, tmp_pxl_out_583, tmp_pxl_out_584, tmp_pxl_out_585, 
tmp_pxl_out_586, tmp_pxl_out_587, tmp_pxl_out_588, tmp_pxl_out_589, tmp_pxl_out_590, tmp_pxl_out_591, tmp_pxl_out_592, tmp_pxl_out_593, tmp_pxl_out_594, 
tmp_pxl_out_595, tmp_pxl_out_596, tmp_pxl_out_597, tmp_pxl_out_598, tmp_pxl_out_599, tmp_pxl_out_600, tmp_pxl_out_601, tmp_pxl_out_602, tmp_pxl_out_603, 
tmp_pxl_out_604, tmp_pxl_out_605, tmp_pxl_out_606, tmp_pxl_out_607, tmp_pxl_out_608, tmp_pxl_out_609, tmp_pxl_out_610, tmp_pxl_out_611, tmp_pxl_out_612, 
tmp_pxl_out_613, tmp_pxl_out_614, tmp_pxl_out_615, tmp_pxl_out_616, tmp_pxl_out_617, tmp_pxl_out_618, tmp_pxl_out_619, tmp_pxl_out_620, tmp_pxl_out_621, 
tmp_pxl_out_622, tmp_pxl_out_623, tmp_pxl_out_624, tmp_pxl_out_625, tmp_pxl_out_626, tmp_pxl_out_627, tmp_pxl_out_628, tmp_pxl_out_629, tmp_pxl_out_630, 
tmp_pxl_out_631, tmp_pxl_out_632, tmp_pxl_out_633, tmp_pxl_out_634, tmp_pxl_out_635, tmp_pxl_out_636, tmp_pxl_out_637, tmp_pxl_out_638, tmp_pxl_out_639, 
tmp_pxl_out_640, tmp_pxl_out_641, tmp_pxl_out_642, tmp_pxl_out_643, tmp_pxl_out_644, tmp_pxl_out_645, tmp_pxl_out_646, tmp_pxl_out_647, tmp_pxl_out_648, 
tmp_pxl_out_649, tmp_pxl_out_650, tmp_pxl_out_651, tmp_pxl_out_652, tmp_pxl_out_653, tmp_pxl_out_654, tmp_pxl_out_655, tmp_pxl_out_656, tmp_pxl_out_657, 
tmp_pxl_out_658, tmp_pxl_out_659, tmp_pxl_out_660, tmp_pxl_out_661, tmp_pxl_out_662, tmp_pxl_out_663, tmp_pxl_out_664, tmp_pxl_out_665, tmp_pxl_out_666, 
tmp_pxl_out_667, tmp_pxl_out_668, tmp_pxl_out_669, tmp_pxl_out_670, tmp_pxl_out_671, tmp_pxl_out_672, tmp_pxl_out_673, tmp_pxl_out_674, tmp_pxl_out_675, 
tmp_pxl_out_676, tmp_pxl_out_677, tmp_pxl_out_678, tmp_pxl_out_679, tmp_pxl_out_680, tmp_pxl_out_681, tmp_pxl_out_682, tmp_pxl_out_683, tmp_pxl_out_684, 
tmp_pxl_out_685, tmp_pxl_out_686, tmp_pxl_out_687, tmp_pxl_out_688, tmp_pxl_out_689, tmp_pxl_out_690, tmp_pxl_out_691, tmp_pxl_out_692, tmp_pxl_out_693, 
tmp_pxl_out_694, tmp_pxl_out_695, tmp_pxl_out_696, tmp_pxl_out_697, tmp_pxl_out_698, tmp_pxl_out_699, tmp_pxl_out_700, tmp_pxl_out_701, tmp_pxl_out_702, 
tmp_pxl_out_703, tmp_pxl_out_704, tmp_pxl_out_705, tmp_pxl_out_706, tmp_pxl_out_707, tmp_pxl_out_708, tmp_pxl_out_709, tmp_pxl_out_710, tmp_pxl_out_711, 
tmp_pxl_out_712, tmp_pxl_out_713, tmp_pxl_out_714, tmp_pxl_out_715, tmp_pxl_out_716, tmp_pxl_out_717, tmp_pxl_out_718, tmp_pxl_out_719, tmp_pxl_out_720, 
tmp_pxl_out_721, tmp_pxl_out_722, tmp_pxl_out_723, tmp_pxl_out_724, tmp_pxl_out_725, tmp_pxl_out_726, tmp_pxl_out_727, tmp_pxl_out_728, tmp_pxl_out_729, 
tmp_pxl_out_730, tmp_pxl_out_731, tmp_pxl_out_732, tmp_pxl_out_733, tmp_pxl_out_734, tmp_pxl_out_735, tmp_pxl_out_736, tmp_pxl_out_737, tmp_pxl_out_738, 
tmp_pxl_out_739, tmp_pxl_out_740, tmp_pxl_out_741, tmp_pxl_out_742, tmp_pxl_out_743, tmp_pxl_out_744, tmp_pxl_out_745, tmp_pxl_out_746, tmp_pxl_out_747, 
tmp_pxl_out_748, tmp_pxl_out_749, tmp_pxl_out_750, tmp_pxl_out_751, tmp_pxl_out_752, tmp_pxl_out_753, tmp_pxl_out_754, tmp_pxl_out_755, tmp_pxl_out_756, 
tmp_pxl_out_757, tmp_pxl_out_758, tmp_pxl_out_759, tmp_pxl_out_760, tmp_pxl_out_761, tmp_pxl_out_762, tmp_pxl_out_763, tmp_pxl_out_764, tmp_pxl_out_765, 
tmp_pxl_out_766, tmp_pxl_out_767, tmp_pxl_out_768, tmp_pxl_out_769, tmp_pxl_out_770, tmp_pxl_out_771, tmp_pxl_out_772, tmp_pxl_out_773, tmp_pxl_out_774, 
tmp_pxl_out_775, tmp_pxl_out_776, tmp_pxl_out_777, tmp_pxl_out_778, tmp_pxl_out_779, tmp_pxl_out_780, tmp_pxl_out_781, tmp_pxl_out_782, tmp_pxl_out_783, 
tmp_pxl_out_784, tmp_pxl_out_785, tmp_pxl_out_786, tmp_pxl_out_787, tmp_pxl_out_788, tmp_pxl_out_789, tmp_pxl_out_790, tmp_pxl_out_791, tmp_pxl_out_792, 
tmp_pxl_out_793, tmp_pxl_out_794, tmp_pxl_out_795, tmp_pxl_out_796, tmp_pxl_out_797, tmp_pxl_out_798, tmp_pxl_out_799, tmp_pxl_out_800, tmp_pxl_out_801, 
tmp_pxl_out_802, tmp_pxl_out_803, tmp_pxl_out_804, tmp_pxl_out_805, tmp_pxl_out_806, tmp_pxl_out_807, tmp_pxl_out_808, tmp_pxl_out_809, tmp_pxl_out_810, 
tmp_pxl_out_811, tmp_pxl_out_812, tmp_pxl_out_813, tmp_pxl_out_814, tmp_pxl_out_815, tmp_pxl_out_816, tmp_pxl_out_817, tmp_pxl_out_818, tmp_pxl_out_819, 
tmp_pxl_out_820, tmp_pxl_out_821, tmp_pxl_out_822, tmp_pxl_out_823, tmp_pxl_out_824, tmp_pxl_out_825, tmp_pxl_out_826, tmp_pxl_out_827, tmp_pxl_out_828, 
tmp_pxl_out_829, tmp_pxl_out_830, tmp_pxl_out_831, tmp_pxl_out_832, tmp_pxl_out_833, tmp_pxl_out_834, tmp_pxl_out_835, tmp_pxl_out_836, tmp_pxl_out_837, 
tmp_pxl_out_838, tmp_pxl_out_839, tmp_pxl_out_840, tmp_pxl_out_841, tmp_pxl_out_842, tmp_pxl_out_843, tmp_pxl_out_844, tmp_pxl_out_845, tmp_pxl_out_846, 
tmp_pxl_out_847, tmp_pxl_out_848, tmp_pxl_out_849, tmp_pxl_out_850, tmp_pxl_out_851, tmp_pxl_out_852, tmp_pxl_out_853, tmp_pxl_out_854, tmp_pxl_out_855, 
tmp_pxl_out_856, tmp_pxl_out_857, tmp_pxl_out_858, tmp_pxl_out_859, tmp_pxl_out_860, tmp_pxl_out_861, tmp_pxl_out_862, tmp_pxl_out_863, tmp_pxl_out_864, 
tmp_pxl_out_865, tmp_pxl_out_866, tmp_pxl_out_867, tmp_pxl_out_868, tmp_pxl_out_869, tmp_pxl_out_870, tmp_pxl_out_871, tmp_pxl_out_872, tmp_pxl_out_873, 
tmp_pxl_out_874, tmp_pxl_out_875, tmp_pxl_out_876, tmp_pxl_out_877, tmp_pxl_out_878, tmp_pxl_out_879, tmp_pxl_out_880, tmp_pxl_out_881, tmp_pxl_out_882, 
tmp_pxl_out_883, tmp_pxl_out_884, tmp_pxl_out_885, tmp_pxl_out_886, tmp_pxl_out_887, tmp_pxl_out_888, tmp_pxl_out_889, tmp_pxl_out_890, tmp_pxl_out_891, 
tmp_pxl_out_892, tmp_pxl_out_893, tmp_pxl_out_894, tmp_pxl_out_895, tmp_pxl_out_896, tmp_pxl_out_897, tmp_pxl_out_898, tmp_pxl_out_899, tmp_pxl_out_900, 
tmp_pxl_out_901, tmp_pxl_out_902, tmp_pxl_out_903, tmp_pxl_out_904, tmp_pxl_out_905, tmp_pxl_out_906, tmp_pxl_out_907, tmp_pxl_out_908, tmp_pxl_out_909, 
tmp_pxl_out_910, tmp_pxl_out_911, tmp_pxl_out_912, tmp_pxl_out_913, tmp_pxl_out_914, tmp_pxl_out_915, tmp_pxl_out_916, tmp_pxl_out_917, tmp_pxl_out_918, 
tmp_pxl_out_919, tmp_pxl_out_920, tmp_pxl_out_921, tmp_pxl_out_922, tmp_pxl_out_923, tmp_pxl_out_924, tmp_pxl_out_925, tmp_pxl_out_926, tmp_pxl_out_927, 
tmp_pxl_out_928, tmp_pxl_out_929, tmp_pxl_out_930, tmp_pxl_out_931, tmp_pxl_out_932, tmp_pxl_out_933, tmp_pxl_out_934, tmp_pxl_out_935, tmp_pxl_out_936, 
tmp_pxl_out_937, tmp_pxl_out_938, tmp_pxl_out_939, tmp_pxl_out_940, tmp_pxl_out_941, tmp_pxl_out_942, tmp_pxl_out_943, tmp_pxl_out_944, tmp_pxl_out_945, 
tmp_pxl_out_946, tmp_pxl_out_947, tmp_pxl_out_948, tmp_pxl_out_949, tmp_pxl_out_950, tmp_pxl_out_951, tmp_pxl_out_952, tmp_pxl_out_953, tmp_pxl_out_954, 
tmp_pxl_out_955, tmp_pxl_out_956, tmp_pxl_out_957, tmp_pxl_out_958, tmp_pxl_out_959, tmp_pxl_out_960, tmp_pxl_out_961, tmp_pxl_out_962, tmp_pxl_out_963, 
tmp_pxl_out_964, tmp_pxl_out_965, tmp_pxl_out_966, tmp_pxl_out_967, tmp_pxl_out_968, tmp_pxl_out_969, tmp_pxl_out_970, tmp_pxl_out_971, tmp_pxl_out_972, 
tmp_pxl_out_973, tmp_pxl_out_974, tmp_pxl_out_975, tmp_pxl_out_976, tmp_pxl_out_977, tmp_pxl_out_978, tmp_pxl_out_979, tmp_pxl_out_980, tmp_pxl_out_981, 
tmp_pxl_out_982, tmp_pxl_out_983, tmp_pxl_out_984, tmp_pxl_out_985, tmp_pxl_out_986, tmp_pxl_out_987, tmp_pxl_out_988, tmp_pxl_out_989, tmp_pxl_out_990, 
tmp_pxl_out_991, tmp_pxl_out_992, tmp_pxl_out_993, tmp_pxl_out_994, tmp_pxl_out_995, tmp_pxl_out_996, tmp_pxl_out_997, tmp_pxl_out_998, tmp_pxl_out_999, 
tmp_pxl_out_1000, tmp_pxl_out_1001, tmp_pxl_out_1002, tmp_pxl_out_1003, tmp_pxl_out_1004, tmp_pxl_out_1005, tmp_pxl_out_1006, tmp_pxl_out_1007, tmp_pxl_out_1008, 
tmp_pxl_out_1009, tmp_pxl_out_1010, tmp_pxl_out_1011, tmp_pxl_out_1012, tmp_pxl_out_1013, tmp_pxl_out_1014, tmp_pxl_out_1015, tmp_pxl_out_1016, tmp_pxl_out_1017, 
tmp_pxl_out_1018, tmp_pxl_out_1019, tmp_pxl_out_1020, tmp_pxl_out_1021, tmp_pxl_out_1022, tmp_pxl_out_1023, tmp_pxl_out_1024;

wire tmp_valid_out_1, tmp_valid_out_2, tmp_valid_out_3, tmp_valid_out_4, tmp_valid_out_5, tmp_valid_out_6, tmp_valid_out_7, tmp_valid_out_8, tmp_valid_out_9, 
tmp_valid_out_10, tmp_valid_out_11, tmp_valid_out_12, tmp_valid_out_13, tmp_valid_out_14, tmp_valid_out_15, tmp_valid_out_16, tmp_valid_out_17, tmp_valid_out_18, 
tmp_valid_out_19, tmp_valid_out_20, tmp_valid_out_21, tmp_valid_out_22, tmp_valid_out_23, tmp_valid_out_24, tmp_valid_out_25, tmp_valid_out_26, tmp_valid_out_27, 
tmp_valid_out_28, tmp_valid_out_29, tmp_valid_out_30, tmp_valid_out_31, tmp_valid_out_32, tmp_valid_out_33, tmp_valid_out_34, tmp_valid_out_35, tmp_valid_out_36, 
tmp_valid_out_37, tmp_valid_out_38, tmp_valid_out_39, tmp_valid_out_40, tmp_valid_out_41, tmp_valid_out_42, tmp_valid_out_43, tmp_valid_out_44, tmp_valid_out_45, 
tmp_valid_out_46, tmp_valid_out_47, tmp_valid_out_48, tmp_valid_out_49, tmp_valid_out_50, tmp_valid_out_51, tmp_valid_out_52, tmp_valid_out_53, tmp_valid_out_54, 
tmp_valid_out_55, tmp_valid_out_56, tmp_valid_out_57, tmp_valid_out_58, tmp_valid_out_59, tmp_valid_out_60, tmp_valid_out_61, tmp_valid_out_62, tmp_valid_out_63, 
tmp_valid_out_64, tmp_valid_out_65, tmp_valid_out_66, tmp_valid_out_67, tmp_valid_out_68, tmp_valid_out_69, tmp_valid_out_70, tmp_valid_out_71, tmp_valid_out_72, 
tmp_valid_out_73, tmp_valid_out_74, tmp_valid_out_75, tmp_valid_out_76, tmp_valid_out_77, tmp_valid_out_78, tmp_valid_out_79, tmp_valid_out_80, tmp_valid_out_81, 
tmp_valid_out_82, tmp_valid_out_83, tmp_valid_out_84, tmp_valid_out_85, tmp_valid_out_86, tmp_valid_out_87, tmp_valid_out_88, tmp_valid_out_89, tmp_valid_out_90, 
tmp_valid_out_91, tmp_valid_out_92, tmp_valid_out_93, tmp_valid_out_94, tmp_valid_out_95, tmp_valid_out_96, tmp_valid_out_97, tmp_valid_out_98, tmp_valid_out_99, 
tmp_valid_out_100, tmp_valid_out_101, tmp_valid_out_102, tmp_valid_out_103, tmp_valid_out_104, tmp_valid_out_105, tmp_valid_out_106, tmp_valid_out_107, tmp_valid_out_108, 
tmp_valid_out_109, tmp_valid_out_110, tmp_valid_out_111, tmp_valid_out_112, tmp_valid_out_113, tmp_valid_out_114, tmp_valid_out_115, tmp_valid_out_116, tmp_valid_out_117, 
tmp_valid_out_118, tmp_valid_out_119, tmp_valid_out_120, tmp_valid_out_121, tmp_valid_out_122, tmp_valid_out_123, tmp_valid_out_124, tmp_valid_out_125, tmp_valid_out_126, 
tmp_valid_out_127, tmp_valid_out_128, tmp_valid_out_129, tmp_valid_out_130, tmp_valid_out_131, tmp_valid_out_132, tmp_valid_out_133, tmp_valid_out_134, tmp_valid_out_135, 
tmp_valid_out_136, tmp_valid_out_137, tmp_valid_out_138, tmp_valid_out_139, tmp_valid_out_140, tmp_valid_out_141, tmp_valid_out_142, tmp_valid_out_143, tmp_valid_out_144, 
tmp_valid_out_145, tmp_valid_out_146, tmp_valid_out_147, tmp_valid_out_148, tmp_valid_out_149, tmp_valid_out_150, tmp_valid_out_151, tmp_valid_out_152, tmp_valid_out_153, 
tmp_valid_out_154, tmp_valid_out_155, tmp_valid_out_156, tmp_valid_out_157, tmp_valid_out_158, tmp_valid_out_159, tmp_valid_out_160, tmp_valid_out_161, tmp_valid_out_162, 
tmp_valid_out_163, tmp_valid_out_164, tmp_valid_out_165, tmp_valid_out_166, tmp_valid_out_167, tmp_valid_out_168, tmp_valid_out_169, tmp_valid_out_170, tmp_valid_out_171, 
tmp_valid_out_172, tmp_valid_out_173, tmp_valid_out_174, tmp_valid_out_175, tmp_valid_out_176, tmp_valid_out_177, tmp_valid_out_178, tmp_valid_out_179, tmp_valid_out_180, 
tmp_valid_out_181, tmp_valid_out_182, tmp_valid_out_183, tmp_valid_out_184, tmp_valid_out_185, tmp_valid_out_186, tmp_valid_out_187, tmp_valid_out_188, tmp_valid_out_189, 
tmp_valid_out_190, tmp_valid_out_191, tmp_valid_out_192, tmp_valid_out_193, tmp_valid_out_194, tmp_valid_out_195, tmp_valid_out_196, tmp_valid_out_197, tmp_valid_out_198, 
tmp_valid_out_199, tmp_valid_out_200, tmp_valid_out_201, tmp_valid_out_202, tmp_valid_out_203, tmp_valid_out_204, tmp_valid_out_205, tmp_valid_out_206, tmp_valid_out_207, 
tmp_valid_out_208, tmp_valid_out_209, tmp_valid_out_210, tmp_valid_out_211, tmp_valid_out_212, tmp_valid_out_213, tmp_valid_out_214, tmp_valid_out_215, tmp_valid_out_216, 
tmp_valid_out_217, tmp_valid_out_218, tmp_valid_out_219, tmp_valid_out_220, tmp_valid_out_221, tmp_valid_out_222, tmp_valid_out_223, tmp_valid_out_224, tmp_valid_out_225, 
tmp_valid_out_226, tmp_valid_out_227, tmp_valid_out_228, tmp_valid_out_229, tmp_valid_out_230, tmp_valid_out_231, tmp_valid_out_232, tmp_valid_out_233, tmp_valid_out_234, 
tmp_valid_out_235, tmp_valid_out_236, tmp_valid_out_237, tmp_valid_out_238, tmp_valid_out_239, tmp_valid_out_240, tmp_valid_out_241, tmp_valid_out_242, tmp_valid_out_243, 
tmp_valid_out_244, tmp_valid_out_245, tmp_valid_out_246, tmp_valid_out_247, tmp_valid_out_248, tmp_valid_out_249, tmp_valid_out_250, tmp_valid_out_251, tmp_valid_out_252, 
tmp_valid_out_253, tmp_valid_out_254, tmp_valid_out_255, tmp_valid_out_256, tmp_valid_out_257, tmp_valid_out_258, tmp_valid_out_259, tmp_valid_out_260, tmp_valid_out_261, 
tmp_valid_out_262, tmp_valid_out_263, tmp_valid_out_264, tmp_valid_out_265, tmp_valid_out_266, tmp_valid_out_267, tmp_valid_out_268, tmp_valid_out_269, tmp_valid_out_270, 
tmp_valid_out_271, tmp_valid_out_272, tmp_valid_out_273, tmp_valid_out_274, tmp_valid_out_275, tmp_valid_out_276, tmp_valid_out_277, tmp_valid_out_278, tmp_valid_out_279, 
tmp_valid_out_280, tmp_valid_out_281, tmp_valid_out_282, tmp_valid_out_283, tmp_valid_out_284, tmp_valid_out_285, tmp_valid_out_286, tmp_valid_out_287, tmp_valid_out_288, 
tmp_valid_out_289, tmp_valid_out_290, tmp_valid_out_291, tmp_valid_out_292, tmp_valid_out_293, tmp_valid_out_294, tmp_valid_out_295, tmp_valid_out_296, tmp_valid_out_297, 
tmp_valid_out_298, tmp_valid_out_299, tmp_valid_out_300, tmp_valid_out_301, tmp_valid_out_302, tmp_valid_out_303, tmp_valid_out_304, tmp_valid_out_305, tmp_valid_out_306, 
tmp_valid_out_307, tmp_valid_out_308, tmp_valid_out_309, tmp_valid_out_310, tmp_valid_out_311, tmp_valid_out_312, tmp_valid_out_313, tmp_valid_out_314, tmp_valid_out_315, 
tmp_valid_out_316, tmp_valid_out_317, tmp_valid_out_318, tmp_valid_out_319, tmp_valid_out_320, tmp_valid_out_321, tmp_valid_out_322, tmp_valid_out_323, tmp_valid_out_324, 
tmp_valid_out_325, tmp_valid_out_326, tmp_valid_out_327, tmp_valid_out_328, tmp_valid_out_329, tmp_valid_out_330, tmp_valid_out_331, tmp_valid_out_332, tmp_valid_out_333, 
tmp_valid_out_334, tmp_valid_out_335, tmp_valid_out_336, tmp_valid_out_337, tmp_valid_out_338, tmp_valid_out_339, tmp_valid_out_340, tmp_valid_out_341, tmp_valid_out_342, 
tmp_valid_out_343, tmp_valid_out_344, tmp_valid_out_345, tmp_valid_out_346, tmp_valid_out_347, tmp_valid_out_348, tmp_valid_out_349, tmp_valid_out_350, tmp_valid_out_351, 
tmp_valid_out_352, tmp_valid_out_353, tmp_valid_out_354, tmp_valid_out_355, tmp_valid_out_356, tmp_valid_out_357, tmp_valid_out_358, tmp_valid_out_359, tmp_valid_out_360, 
tmp_valid_out_361, tmp_valid_out_362, tmp_valid_out_363, tmp_valid_out_364, tmp_valid_out_365, tmp_valid_out_366, tmp_valid_out_367, tmp_valid_out_368, tmp_valid_out_369, 
tmp_valid_out_370, tmp_valid_out_371, tmp_valid_out_372, tmp_valid_out_373, tmp_valid_out_374, tmp_valid_out_375, tmp_valid_out_376, tmp_valid_out_377, tmp_valid_out_378, 
tmp_valid_out_379, tmp_valid_out_380, tmp_valid_out_381, tmp_valid_out_382, tmp_valid_out_383, tmp_valid_out_384, tmp_valid_out_385, tmp_valid_out_386, tmp_valid_out_387, 
tmp_valid_out_388, tmp_valid_out_389, tmp_valid_out_390, tmp_valid_out_391, tmp_valid_out_392, tmp_valid_out_393, tmp_valid_out_394, tmp_valid_out_395, tmp_valid_out_396, 
tmp_valid_out_397, tmp_valid_out_398, tmp_valid_out_399, tmp_valid_out_400, tmp_valid_out_401, tmp_valid_out_402, tmp_valid_out_403, tmp_valid_out_404, tmp_valid_out_405, 
tmp_valid_out_406, tmp_valid_out_407, tmp_valid_out_408, tmp_valid_out_409, tmp_valid_out_410, tmp_valid_out_411, tmp_valid_out_412, tmp_valid_out_413, tmp_valid_out_414, 
tmp_valid_out_415, tmp_valid_out_416, tmp_valid_out_417, tmp_valid_out_418, tmp_valid_out_419, tmp_valid_out_420, tmp_valid_out_421, tmp_valid_out_422, tmp_valid_out_423, 
tmp_valid_out_424, tmp_valid_out_425, tmp_valid_out_426, tmp_valid_out_427, tmp_valid_out_428, tmp_valid_out_429, tmp_valid_out_430, tmp_valid_out_431, tmp_valid_out_432, 
tmp_valid_out_433, tmp_valid_out_434, tmp_valid_out_435, tmp_valid_out_436, tmp_valid_out_437, tmp_valid_out_438, tmp_valid_out_439, tmp_valid_out_440, tmp_valid_out_441, 
tmp_valid_out_442, tmp_valid_out_443, tmp_valid_out_444, tmp_valid_out_445, tmp_valid_out_446, tmp_valid_out_447, tmp_valid_out_448, tmp_valid_out_449, tmp_valid_out_450, 
tmp_valid_out_451, tmp_valid_out_452, tmp_valid_out_453, tmp_valid_out_454, tmp_valid_out_455, tmp_valid_out_456, tmp_valid_out_457, tmp_valid_out_458, tmp_valid_out_459, 
tmp_valid_out_460, tmp_valid_out_461, tmp_valid_out_462, tmp_valid_out_463, tmp_valid_out_464, tmp_valid_out_465, tmp_valid_out_466, tmp_valid_out_467, tmp_valid_out_468, 
tmp_valid_out_469, tmp_valid_out_470, tmp_valid_out_471, tmp_valid_out_472, tmp_valid_out_473, tmp_valid_out_474, tmp_valid_out_475, tmp_valid_out_476, tmp_valid_out_477, 
tmp_valid_out_478, tmp_valid_out_479, tmp_valid_out_480, tmp_valid_out_481, tmp_valid_out_482, tmp_valid_out_483, tmp_valid_out_484, tmp_valid_out_485, tmp_valid_out_486, 
tmp_valid_out_487, tmp_valid_out_488, tmp_valid_out_489, tmp_valid_out_490, tmp_valid_out_491, tmp_valid_out_492, tmp_valid_out_493, tmp_valid_out_494, tmp_valid_out_495, 
tmp_valid_out_496, tmp_valid_out_497, tmp_valid_out_498, tmp_valid_out_499, tmp_valid_out_500, tmp_valid_out_501, tmp_valid_out_502, tmp_valid_out_503, tmp_valid_out_504, 
tmp_valid_out_505, tmp_valid_out_506, tmp_valid_out_507, tmp_valid_out_508, tmp_valid_out_509, tmp_valid_out_510, tmp_valid_out_511, tmp_valid_out_512, tmp_valid_out_513, 
tmp_valid_out_514, tmp_valid_out_515, tmp_valid_out_516, tmp_valid_out_517, tmp_valid_out_518, tmp_valid_out_519, tmp_valid_out_520, tmp_valid_out_521, tmp_valid_out_522, 
tmp_valid_out_523, tmp_valid_out_524, tmp_valid_out_525, tmp_valid_out_526, tmp_valid_out_527, tmp_valid_out_528, tmp_valid_out_529, tmp_valid_out_530, tmp_valid_out_531, 
tmp_valid_out_532, tmp_valid_out_533, tmp_valid_out_534, tmp_valid_out_535, tmp_valid_out_536, tmp_valid_out_537, tmp_valid_out_538, tmp_valid_out_539, tmp_valid_out_540, 
tmp_valid_out_541, tmp_valid_out_542, tmp_valid_out_543, tmp_valid_out_544, tmp_valid_out_545, tmp_valid_out_546, tmp_valid_out_547, tmp_valid_out_548, tmp_valid_out_549, 
tmp_valid_out_550, tmp_valid_out_551, tmp_valid_out_552, tmp_valid_out_553, tmp_valid_out_554, tmp_valid_out_555, tmp_valid_out_556, tmp_valid_out_557, tmp_valid_out_558, 
tmp_valid_out_559, tmp_valid_out_560, tmp_valid_out_561, tmp_valid_out_562, tmp_valid_out_563, tmp_valid_out_564, tmp_valid_out_565, tmp_valid_out_566, tmp_valid_out_567, 
tmp_valid_out_568, tmp_valid_out_569, tmp_valid_out_570, tmp_valid_out_571, tmp_valid_out_572, tmp_valid_out_573, tmp_valid_out_574, tmp_valid_out_575, tmp_valid_out_576, 
tmp_valid_out_577, tmp_valid_out_578, tmp_valid_out_579, tmp_valid_out_580, tmp_valid_out_581, tmp_valid_out_582, tmp_valid_out_583, tmp_valid_out_584, tmp_valid_out_585, 
tmp_valid_out_586, tmp_valid_out_587, tmp_valid_out_588, tmp_valid_out_589, tmp_valid_out_590, tmp_valid_out_591, tmp_valid_out_592, tmp_valid_out_593, tmp_valid_out_594, 
tmp_valid_out_595, tmp_valid_out_596, tmp_valid_out_597, tmp_valid_out_598, tmp_valid_out_599, tmp_valid_out_600, tmp_valid_out_601, tmp_valid_out_602, tmp_valid_out_603, 
tmp_valid_out_604, tmp_valid_out_605, tmp_valid_out_606, tmp_valid_out_607, tmp_valid_out_608, tmp_valid_out_609, tmp_valid_out_610, tmp_valid_out_611, tmp_valid_out_612, 
tmp_valid_out_613, tmp_valid_out_614, tmp_valid_out_615, tmp_valid_out_616, tmp_valid_out_617, tmp_valid_out_618, tmp_valid_out_619, tmp_valid_out_620, tmp_valid_out_621, 
tmp_valid_out_622, tmp_valid_out_623, tmp_valid_out_624, tmp_valid_out_625, tmp_valid_out_626, tmp_valid_out_627, tmp_valid_out_628, tmp_valid_out_629, tmp_valid_out_630, 
tmp_valid_out_631, tmp_valid_out_632, tmp_valid_out_633, tmp_valid_out_634, tmp_valid_out_635, tmp_valid_out_636, tmp_valid_out_637, tmp_valid_out_638, tmp_valid_out_639, 
tmp_valid_out_640, tmp_valid_out_641, tmp_valid_out_642, tmp_valid_out_643, tmp_valid_out_644, tmp_valid_out_645, tmp_valid_out_646, tmp_valid_out_647, tmp_valid_out_648, 
tmp_valid_out_649, tmp_valid_out_650, tmp_valid_out_651, tmp_valid_out_652, tmp_valid_out_653, tmp_valid_out_654, tmp_valid_out_655, tmp_valid_out_656, tmp_valid_out_657, 
tmp_valid_out_658, tmp_valid_out_659, tmp_valid_out_660, tmp_valid_out_661, tmp_valid_out_662, tmp_valid_out_663, tmp_valid_out_664, tmp_valid_out_665, tmp_valid_out_666, 
tmp_valid_out_667, tmp_valid_out_668, tmp_valid_out_669, tmp_valid_out_670, tmp_valid_out_671, tmp_valid_out_672, tmp_valid_out_673, tmp_valid_out_674, tmp_valid_out_675, 
tmp_valid_out_676, tmp_valid_out_677, tmp_valid_out_678, tmp_valid_out_679, tmp_valid_out_680, tmp_valid_out_681, tmp_valid_out_682, tmp_valid_out_683, tmp_valid_out_684, 
tmp_valid_out_685, tmp_valid_out_686, tmp_valid_out_687, tmp_valid_out_688, tmp_valid_out_689, tmp_valid_out_690, tmp_valid_out_691, tmp_valid_out_692, tmp_valid_out_693, 
tmp_valid_out_694, tmp_valid_out_695, tmp_valid_out_696, tmp_valid_out_697, tmp_valid_out_698, tmp_valid_out_699, tmp_valid_out_700, tmp_valid_out_701, tmp_valid_out_702, 
tmp_valid_out_703, tmp_valid_out_704, tmp_valid_out_705, tmp_valid_out_706, tmp_valid_out_707, tmp_valid_out_708, tmp_valid_out_709, tmp_valid_out_710, tmp_valid_out_711, 
tmp_valid_out_712, tmp_valid_out_713, tmp_valid_out_714, tmp_valid_out_715, tmp_valid_out_716, tmp_valid_out_717, tmp_valid_out_718, tmp_valid_out_719, tmp_valid_out_720, 
tmp_valid_out_721, tmp_valid_out_722, tmp_valid_out_723, tmp_valid_out_724, tmp_valid_out_725, tmp_valid_out_726, tmp_valid_out_727, tmp_valid_out_728, tmp_valid_out_729, 
tmp_valid_out_730, tmp_valid_out_731, tmp_valid_out_732, tmp_valid_out_733, tmp_valid_out_734, tmp_valid_out_735, tmp_valid_out_736, tmp_valid_out_737, tmp_valid_out_738, 
tmp_valid_out_739, tmp_valid_out_740, tmp_valid_out_741, tmp_valid_out_742, tmp_valid_out_743, tmp_valid_out_744, tmp_valid_out_745, tmp_valid_out_746, tmp_valid_out_747, 
tmp_valid_out_748, tmp_valid_out_749, tmp_valid_out_750, tmp_valid_out_751, tmp_valid_out_752, tmp_valid_out_753, tmp_valid_out_754, tmp_valid_out_755, tmp_valid_out_756, 
tmp_valid_out_757, tmp_valid_out_758, tmp_valid_out_759, tmp_valid_out_760, tmp_valid_out_761, tmp_valid_out_762, tmp_valid_out_763, tmp_valid_out_764, tmp_valid_out_765, 
tmp_valid_out_766, tmp_valid_out_767, tmp_valid_out_768, tmp_valid_out_769, tmp_valid_out_770, tmp_valid_out_771, tmp_valid_out_772, tmp_valid_out_773, tmp_valid_out_774, 
tmp_valid_out_775, tmp_valid_out_776, tmp_valid_out_777, tmp_valid_out_778, tmp_valid_out_779, tmp_valid_out_780, tmp_valid_out_781, tmp_valid_out_782, tmp_valid_out_783, 
tmp_valid_out_784, tmp_valid_out_785, tmp_valid_out_786, tmp_valid_out_787, tmp_valid_out_788, tmp_valid_out_789, tmp_valid_out_790, tmp_valid_out_791, tmp_valid_out_792, 
tmp_valid_out_793, tmp_valid_out_794, tmp_valid_out_795, tmp_valid_out_796, tmp_valid_out_797, tmp_valid_out_798, tmp_valid_out_799, tmp_valid_out_800, tmp_valid_out_801, 
tmp_valid_out_802, tmp_valid_out_803, tmp_valid_out_804, tmp_valid_out_805, tmp_valid_out_806, tmp_valid_out_807, tmp_valid_out_808, tmp_valid_out_809, tmp_valid_out_810, 
tmp_valid_out_811, tmp_valid_out_812, tmp_valid_out_813, tmp_valid_out_814, tmp_valid_out_815, tmp_valid_out_816, tmp_valid_out_817, tmp_valid_out_818, tmp_valid_out_819, 
tmp_valid_out_820, tmp_valid_out_821, tmp_valid_out_822, tmp_valid_out_823, tmp_valid_out_824, tmp_valid_out_825, tmp_valid_out_826, tmp_valid_out_827, tmp_valid_out_828, 
tmp_valid_out_829, tmp_valid_out_830, tmp_valid_out_831, tmp_valid_out_832, tmp_valid_out_833, tmp_valid_out_834, tmp_valid_out_835, tmp_valid_out_836, tmp_valid_out_837, 
tmp_valid_out_838, tmp_valid_out_839, tmp_valid_out_840, tmp_valid_out_841, tmp_valid_out_842, tmp_valid_out_843, tmp_valid_out_844, tmp_valid_out_845, tmp_valid_out_846, 
tmp_valid_out_847, tmp_valid_out_848, tmp_valid_out_849, tmp_valid_out_850, tmp_valid_out_851, tmp_valid_out_852, tmp_valid_out_853, tmp_valid_out_854, tmp_valid_out_855, 
tmp_valid_out_856, tmp_valid_out_857, tmp_valid_out_858, tmp_valid_out_859, tmp_valid_out_860, tmp_valid_out_861, tmp_valid_out_862, tmp_valid_out_863, tmp_valid_out_864, 
tmp_valid_out_865, tmp_valid_out_866, tmp_valid_out_867, tmp_valid_out_868, tmp_valid_out_869, tmp_valid_out_870, tmp_valid_out_871, tmp_valid_out_872, tmp_valid_out_873, 
tmp_valid_out_874, tmp_valid_out_875, tmp_valid_out_876, tmp_valid_out_877, tmp_valid_out_878, tmp_valid_out_879, tmp_valid_out_880, tmp_valid_out_881, tmp_valid_out_882, 
tmp_valid_out_883, tmp_valid_out_884, tmp_valid_out_885, tmp_valid_out_886, tmp_valid_out_887, tmp_valid_out_888, tmp_valid_out_889, tmp_valid_out_890, tmp_valid_out_891, 
tmp_valid_out_892, tmp_valid_out_893, tmp_valid_out_894, tmp_valid_out_895, tmp_valid_out_896, tmp_valid_out_897, tmp_valid_out_898, tmp_valid_out_899, tmp_valid_out_900, 
tmp_valid_out_901, tmp_valid_out_902, tmp_valid_out_903, tmp_valid_out_904, tmp_valid_out_905, tmp_valid_out_906, tmp_valid_out_907, tmp_valid_out_908, tmp_valid_out_909, 
tmp_valid_out_910, tmp_valid_out_911, tmp_valid_out_912, tmp_valid_out_913, tmp_valid_out_914, tmp_valid_out_915, tmp_valid_out_916, tmp_valid_out_917, tmp_valid_out_918, 
tmp_valid_out_919, tmp_valid_out_920, tmp_valid_out_921, tmp_valid_out_922, tmp_valid_out_923, tmp_valid_out_924, tmp_valid_out_925, tmp_valid_out_926, tmp_valid_out_927, 
tmp_valid_out_928, tmp_valid_out_929, tmp_valid_out_930, tmp_valid_out_931, tmp_valid_out_932, tmp_valid_out_933, tmp_valid_out_934, tmp_valid_out_935, tmp_valid_out_936, 
tmp_valid_out_937, tmp_valid_out_938, tmp_valid_out_939, tmp_valid_out_940, tmp_valid_out_941, tmp_valid_out_942, tmp_valid_out_943, tmp_valid_out_944, tmp_valid_out_945, 
tmp_valid_out_946, tmp_valid_out_947, tmp_valid_out_948, tmp_valid_out_949, tmp_valid_out_950, tmp_valid_out_951, tmp_valid_out_952, tmp_valid_out_953, tmp_valid_out_954, 
tmp_valid_out_955, tmp_valid_out_956, tmp_valid_out_957, tmp_valid_out_958, tmp_valid_out_959, tmp_valid_out_960, tmp_valid_out_961, tmp_valid_out_962, tmp_valid_out_963, 
tmp_valid_out_964, tmp_valid_out_965, tmp_valid_out_966, tmp_valid_out_967, tmp_valid_out_968, tmp_valid_out_969, tmp_valid_out_970, tmp_valid_out_971, tmp_valid_out_972, 
tmp_valid_out_973, tmp_valid_out_974, tmp_valid_out_975, tmp_valid_out_976, tmp_valid_out_977, tmp_valid_out_978, tmp_valid_out_979, tmp_valid_out_980, tmp_valid_out_981, 
tmp_valid_out_982, tmp_valid_out_983, tmp_valid_out_984, tmp_valid_out_985, tmp_valid_out_986, tmp_valid_out_987, tmp_valid_out_988, tmp_valid_out_989, tmp_valid_out_990, 
tmp_valid_out_991, tmp_valid_out_992, tmp_valid_out_993, tmp_valid_out_994, tmp_valid_out_995, tmp_valid_out_996, tmp_valid_out_997, tmp_valid_out_998, tmp_valid_out_999, 
tmp_valid_out_1000, tmp_valid_out_1001, tmp_valid_out_1002, tmp_valid_out_1003, tmp_valid_out_1004, tmp_valid_out_1005, tmp_valid_out_1006, tmp_valid_out_1007, tmp_valid_out_1008, 
tmp_valid_out_1009, tmp_valid_out_1010, tmp_valid_out_1011, tmp_valid_out_1012, tmp_valid_out_1013, tmp_valid_out_1014, tmp_valid_out_1015, tmp_valid_out_1016, tmp_valid_out_1017, 
tmp_valid_out_1018, tmp_valid_out_1019, tmp_valid_out_1020, tmp_valid_out_1021, tmp_valid_out_1022, tmp_valid_out_1023, tmp_valid_out_1024;

Conv2d_2a_3x3_32 #(D,DATA_WIDTH) uut1 (

clk, 
reset, 
valid_in_1,valid_in_2,valid_in_3,valid_in_4,valid_in_5,valid_in_6,valid_in_7,valid_in_8,valid_in_9,
valid_in_10,valid_in_11,valid_in_12,valid_in_13,valid_in_14,valid_in_15,valid_in_16,valid_in_17,valid_in_18,
valid_in_19,valid_in_20,valid_in_21,valid_in_22,valid_in_23,valid_in_24,valid_in_25,valid_in_26,valid_in_27,
valid_in_28,valid_in_29,valid_in_30,valid_in_31,valid_in_32,

pxl_in_1,pxl_in_2,pxl_in_3,pxl_in_4,pxl_in_5,pxl_in_6,pxl_in_7,pxl_in_8,pxl_in_9,
pxl_in_10,pxl_in_11,pxl_in_12,pxl_in_13,pxl_in_14,pxl_in_15,pxl_in_16,pxl_in_17,pxl_in_18,
pxl_in_19,pxl_in_20,pxl_in_21,pxl_in_22,pxl_in_23,pxl_in_24,pxl_in_25,pxl_in_26,pxl_in_27,
pxl_in_28,pxl_in_29,pxl_in_30,pxl_in_31,pxl_in_32,
                             		
tmp_pxl_out_1, tmp_pxl_out_2, tmp_pxl_out_3, tmp_pxl_out_4, tmp_pxl_out_5, tmp_pxl_out_6, tmp_pxl_out_7, tmp_pxl_out_8, tmp_pxl_out_9, 
tmp_pxl_out_10, tmp_pxl_out_11, tmp_pxl_out_12, tmp_pxl_out_13, tmp_pxl_out_14, tmp_pxl_out_15, tmp_pxl_out_16, tmp_pxl_out_17, tmp_pxl_out_18, 
tmp_pxl_out_19, tmp_pxl_out_20, tmp_pxl_out_21, tmp_pxl_out_22, tmp_pxl_out_23, tmp_pxl_out_24, tmp_pxl_out_25, tmp_pxl_out_26, tmp_pxl_out_27, 
tmp_pxl_out_28, tmp_pxl_out_29, tmp_pxl_out_30, tmp_pxl_out_31, tmp_pxl_out_32, tmp_pxl_out_33, tmp_pxl_out_34, tmp_pxl_out_35, tmp_pxl_out_36, 
tmp_pxl_out_37, tmp_pxl_out_38, tmp_pxl_out_39, tmp_pxl_out_40, tmp_pxl_out_41, tmp_pxl_out_42, tmp_pxl_out_43, tmp_pxl_out_44, tmp_pxl_out_45, 
tmp_pxl_out_46, tmp_pxl_out_47, tmp_pxl_out_48, tmp_pxl_out_49, tmp_pxl_out_50, tmp_pxl_out_51, tmp_pxl_out_52, tmp_pxl_out_53, tmp_pxl_out_54, 
tmp_pxl_out_55, tmp_pxl_out_56, tmp_pxl_out_57, tmp_pxl_out_58, tmp_pxl_out_59, tmp_pxl_out_60, tmp_pxl_out_61, tmp_pxl_out_62, tmp_pxl_out_63, 
tmp_pxl_out_64, tmp_pxl_out_65, tmp_pxl_out_66, tmp_pxl_out_67, tmp_pxl_out_68, tmp_pxl_out_69, tmp_pxl_out_70, tmp_pxl_out_71, tmp_pxl_out_72, 
tmp_pxl_out_73, tmp_pxl_out_74, tmp_pxl_out_75, tmp_pxl_out_76, tmp_pxl_out_77, tmp_pxl_out_78, tmp_pxl_out_79, tmp_pxl_out_80, tmp_pxl_out_81, 
tmp_pxl_out_82, tmp_pxl_out_83, tmp_pxl_out_84, tmp_pxl_out_85, tmp_pxl_out_86, tmp_pxl_out_87, tmp_pxl_out_88, tmp_pxl_out_89, tmp_pxl_out_90, 
tmp_pxl_out_91, tmp_pxl_out_92, tmp_pxl_out_93, tmp_pxl_out_94, tmp_pxl_out_95, tmp_pxl_out_96, tmp_pxl_out_97, tmp_pxl_out_98, tmp_pxl_out_99, 
tmp_pxl_out_100, tmp_pxl_out_101, tmp_pxl_out_102, tmp_pxl_out_103, tmp_pxl_out_104, tmp_pxl_out_105, tmp_pxl_out_106, tmp_pxl_out_107, tmp_pxl_out_108, 
tmp_pxl_out_109, tmp_pxl_out_110, tmp_pxl_out_111, tmp_pxl_out_112, tmp_pxl_out_113, tmp_pxl_out_114, tmp_pxl_out_115, tmp_pxl_out_116, tmp_pxl_out_117, 
tmp_pxl_out_118, tmp_pxl_out_119, tmp_pxl_out_120, tmp_pxl_out_121, tmp_pxl_out_122, tmp_pxl_out_123, tmp_pxl_out_124, tmp_pxl_out_125, tmp_pxl_out_126, 
tmp_pxl_out_127, tmp_pxl_out_128, tmp_pxl_out_129, tmp_pxl_out_130, tmp_pxl_out_131, tmp_pxl_out_132, tmp_pxl_out_133, tmp_pxl_out_134, tmp_pxl_out_135, 
tmp_pxl_out_136, tmp_pxl_out_137, tmp_pxl_out_138, tmp_pxl_out_139, tmp_pxl_out_140, tmp_pxl_out_141, tmp_pxl_out_142, tmp_pxl_out_143, tmp_pxl_out_144, 
tmp_pxl_out_145, tmp_pxl_out_146, tmp_pxl_out_147, tmp_pxl_out_148, tmp_pxl_out_149, tmp_pxl_out_150, tmp_pxl_out_151, tmp_pxl_out_152, tmp_pxl_out_153, 
tmp_pxl_out_154, tmp_pxl_out_155, tmp_pxl_out_156, tmp_pxl_out_157, tmp_pxl_out_158, tmp_pxl_out_159, tmp_pxl_out_160, tmp_pxl_out_161, tmp_pxl_out_162, 
tmp_pxl_out_163, tmp_pxl_out_164, tmp_pxl_out_165, tmp_pxl_out_166, tmp_pxl_out_167, tmp_pxl_out_168, tmp_pxl_out_169, tmp_pxl_out_170, tmp_pxl_out_171, 
tmp_pxl_out_172, tmp_pxl_out_173, tmp_pxl_out_174, tmp_pxl_out_175, tmp_pxl_out_176, tmp_pxl_out_177, tmp_pxl_out_178, tmp_pxl_out_179, tmp_pxl_out_180, 
tmp_pxl_out_181, tmp_pxl_out_182, tmp_pxl_out_183, tmp_pxl_out_184, tmp_pxl_out_185, tmp_pxl_out_186, tmp_pxl_out_187, tmp_pxl_out_188, tmp_pxl_out_189, 
tmp_pxl_out_190, tmp_pxl_out_191, tmp_pxl_out_192, tmp_pxl_out_193, tmp_pxl_out_194, tmp_pxl_out_195, tmp_pxl_out_196, tmp_pxl_out_197, tmp_pxl_out_198, 
tmp_pxl_out_199, tmp_pxl_out_200, tmp_pxl_out_201, tmp_pxl_out_202, tmp_pxl_out_203, tmp_pxl_out_204, tmp_pxl_out_205, tmp_pxl_out_206, tmp_pxl_out_207, 
tmp_pxl_out_208, tmp_pxl_out_209, tmp_pxl_out_210, tmp_pxl_out_211, tmp_pxl_out_212, tmp_pxl_out_213, tmp_pxl_out_214, tmp_pxl_out_215, tmp_pxl_out_216, 
tmp_pxl_out_217, tmp_pxl_out_218, tmp_pxl_out_219, tmp_pxl_out_220, tmp_pxl_out_221, tmp_pxl_out_222, tmp_pxl_out_223, tmp_pxl_out_224, tmp_pxl_out_225, 
tmp_pxl_out_226, tmp_pxl_out_227, tmp_pxl_out_228, tmp_pxl_out_229, tmp_pxl_out_230, tmp_pxl_out_231, tmp_pxl_out_232, tmp_pxl_out_233, tmp_pxl_out_234, 
tmp_pxl_out_235, tmp_pxl_out_236, tmp_pxl_out_237, tmp_pxl_out_238, tmp_pxl_out_239, tmp_pxl_out_240, tmp_pxl_out_241, tmp_pxl_out_242, tmp_pxl_out_243, 
tmp_pxl_out_244, tmp_pxl_out_245, tmp_pxl_out_246, tmp_pxl_out_247, tmp_pxl_out_248, tmp_pxl_out_249, tmp_pxl_out_250, tmp_pxl_out_251, tmp_pxl_out_252, 
tmp_pxl_out_253, tmp_pxl_out_254, tmp_pxl_out_255, tmp_pxl_out_256, tmp_pxl_out_257, tmp_pxl_out_258, tmp_pxl_out_259, tmp_pxl_out_260, tmp_pxl_out_261, 
tmp_pxl_out_262, tmp_pxl_out_263, tmp_pxl_out_264, tmp_pxl_out_265, tmp_pxl_out_266, tmp_pxl_out_267, tmp_pxl_out_268, tmp_pxl_out_269, tmp_pxl_out_270, 
tmp_pxl_out_271, tmp_pxl_out_272, tmp_pxl_out_273, tmp_pxl_out_274, tmp_pxl_out_275, tmp_pxl_out_276, tmp_pxl_out_277, tmp_pxl_out_278, tmp_pxl_out_279, 
tmp_pxl_out_280, tmp_pxl_out_281, tmp_pxl_out_282, tmp_pxl_out_283, tmp_pxl_out_284, tmp_pxl_out_285, tmp_pxl_out_286, tmp_pxl_out_287, tmp_pxl_out_288, 
tmp_pxl_out_289, tmp_pxl_out_290, tmp_pxl_out_291, tmp_pxl_out_292, tmp_pxl_out_293, tmp_pxl_out_294, tmp_pxl_out_295, tmp_pxl_out_296, tmp_pxl_out_297, 
tmp_pxl_out_298, tmp_pxl_out_299, tmp_pxl_out_300, tmp_pxl_out_301, tmp_pxl_out_302, tmp_pxl_out_303, tmp_pxl_out_304, tmp_pxl_out_305, tmp_pxl_out_306, 
tmp_pxl_out_307, tmp_pxl_out_308, tmp_pxl_out_309, tmp_pxl_out_310, tmp_pxl_out_311, tmp_pxl_out_312, tmp_pxl_out_313, tmp_pxl_out_314, tmp_pxl_out_315, 
tmp_pxl_out_316, tmp_pxl_out_317, tmp_pxl_out_318, tmp_pxl_out_319, tmp_pxl_out_320, tmp_pxl_out_321, tmp_pxl_out_322, tmp_pxl_out_323, tmp_pxl_out_324, 
tmp_pxl_out_325, tmp_pxl_out_326, tmp_pxl_out_327, tmp_pxl_out_328, tmp_pxl_out_329, tmp_pxl_out_330, tmp_pxl_out_331, tmp_pxl_out_332, tmp_pxl_out_333, 
tmp_pxl_out_334, tmp_pxl_out_335, tmp_pxl_out_336, tmp_pxl_out_337, tmp_pxl_out_338, tmp_pxl_out_339, tmp_pxl_out_340, tmp_pxl_out_341, tmp_pxl_out_342, 
tmp_pxl_out_343, tmp_pxl_out_344, tmp_pxl_out_345, tmp_pxl_out_346, tmp_pxl_out_347, tmp_pxl_out_348, tmp_pxl_out_349, tmp_pxl_out_350, tmp_pxl_out_351, 
tmp_pxl_out_352, tmp_pxl_out_353, tmp_pxl_out_354, tmp_pxl_out_355, tmp_pxl_out_356, tmp_pxl_out_357, tmp_pxl_out_358, tmp_pxl_out_359, tmp_pxl_out_360, 
tmp_pxl_out_361, tmp_pxl_out_362, tmp_pxl_out_363, tmp_pxl_out_364, tmp_pxl_out_365, tmp_pxl_out_366, tmp_pxl_out_367, tmp_pxl_out_368, tmp_pxl_out_369, 
tmp_pxl_out_370, tmp_pxl_out_371, tmp_pxl_out_372, tmp_pxl_out_373, tmp_pxl_out_374, tmp_pxl_out_375, tmp_pxl_out_376, tmp_pxl_out_377, tmp_pxl_out_378, 
tmp_pxl_out_379, tmp_pxl_out_380, tmp_pxl_out_381, tmp_pxl_out_382, tmp_pxl_out_383, tmp_pxl_out_384, tmp_pxl_out_385, tmp_pxl_out_386, tmp_pxl_out_387, 
tmp_pxl_out_388, tmp_pxl_out_389, tmp_pxl_out_390, tmp_pxl_out_391, tmp_pxl_out_392, tmp_pxl_out_393, tmp_pxl_out_394, tmp_pxl_out_395, tmp_pxl_out_396, 
tmp_pxl_out_397, tmp_pxl_out_398, tmp_pxl_out_399, tmp_pxl_out_400, tmp_pxl_out_401, tmp_pxl_out_402, tmp_pxl_out_403, tmp_pxl_out_404, tmp_pxl_out_405, 
tmp_pxl_out_406, tmp_pxl_out_407, tmp_pxl_out_408, tmp_pxl_out_409, tmp_pxl_out_410, tmp_pxl_out_411, tmp_pxl_out_412, tmp_pxl_out_413, tmp_pxl_out_414, 
tmp_pxl_out_415, tmp_pxl_out_416, tmp_pxl_out_417, tmp_pxl_out_418, tmp_pxl_out_419, tmp_pxl_out_420, tmp_pxl_out_421, tmp_pxl_out_422, tmp_pxl_out_423, 
tmp_pxl_out_424, tmp_pxl_out_425, tmp_pxl_out_426, tmp_pxl_out_427, tmp_pxl_out_428, tmp_pxl_out_429, tmp_pxl_out_430, tmp_pxl_out_431, tmp_pxl_out_432, 
tmp_pxl_out_433, tmp_pxl_out_434, tmp_pxl_out_435, tmp_pxl_out_436, tmp_pxl_out_437, tmp_pxl_out_438, tmp_pxl_out_439, tmp_pxl_out_440, tmp_pxl_out_441, 
tmp_pxl_out_442, tmp_pxl_out_443, tmp_pxl_out_444, tmp_pxl_out_445, tmp_pxl_out_446, tmp_pxl_out_447, tmp_pxl_out_448, tmp_pxl_out_449, tmp_pxl_out_450, 
tmp_pxl_out_451, tmp_pxl_out_452, tmp_pxl_out_453, tmp_pxl_out_454, tmp_pxl_out_455, tmp_pxl_out_456, tmp_pxl_out_457, tmp_pxl_out_458, tmp_pxl_out_459, 
tmp_pxl_out_460, tmp_pxl_out_461, tmp_pxl_out_462, tmp_pxl_out_463, tmp_pxl_out_464, tmp_pxl_out_465, tmp_pxl_out_466, tmp_pxl_out_467, tmp_pxl_out_468, 
tmp_pxl_out_469, tmp_pxl_out_470, tmp_pxl_out_471, tmp_pxl_out_472, tmp_pxl_out_473, tmp_pxl_out_474, tmp_pxl_out_475, tmp_pxl_out_476, tmp_pxl_out_477, 
tmp_pxl_out_478, tmp_pxl_out_479, tmp_pxl_out_480, tmp_pxl_out_481, tmp_pxl_out_482, tmp_pxl_out_483, tmp_pxl_out_484, tmp_pxl_out_485, tmp_pxl_out_486, 
tmp_pxl_out_487, tmp_pxl_out_488, tmp_pxl_out_489, tmp_pxl_out_490, tmp_pxl_out_491, tmp_pxl_out_492, tmp_pxl_out_493, tmp_pxl_out_494, tmp_pxl_out_495, 
tmp_pxl_out_496, tmp_pxl_out_497, tmp_pxl_out_498, tmp_pxl_out_499, tmp_pxl_out_500, tmp_pxl_out_501, tmp_pxl_out_502, tmp_pxl_out_503, tmp_pxl_out_504, 
tmp_pxl_out_505, tmp_pxl_out_506, tmp_pxl_out_507, tmp_pxl_out_508, tmp_pxl_out_509, tmp_pxl_out_510, tmp_pxl_out_511, tmp_pxl_out_512, tmp_pxl_out_513, 
tmp_pxl_out_514, tmp_pxl_out_515, tmp_pxl_out_516, tmp_pxl_out_517, tmp_pxl_out_518, tmp_pxl_out_519, tmp_pxl_out_520, tmp_pxl_out_521, tmp_pxl_out_522, 
tmp_pxl_out_523, tmp_pxl_out_524, tmp_pxl_out_525, tmp_pxl_out_526, tmp_pxl_out_527, tmp_pxl_out_528, tmp_pxl_out_529, tmp_pxl_out_530, tmp_pxl_out_531, 
tmp_pxl_out_532, tmp_pxl_out_533, tmp_pxl_out_534, tmp_pxl_out_535, tmp_pxl_out_536, tmp_pxl_out_537, tmp_pxl_out_538, tmp_pxl_out_539, tmp_pxl_out_540, 
tmp_pxl_out_541, tmp_pxl_out_542, tmp_pxl_out_543, tmp_pxl_out_544, tmp_pxl_out_545, tmp_pxl_out_546, tmp_pxl_out_547, tmp_pxl_out_548, tmp_pxl_out_549, 
tmp_pxl_out_550, tmp_pxl_out_551, tmp_pxl_out_552, tmp_pxl_out_553, tmp_pxl_out_554, tmp_pxl_out_555, tmp_pxl_out_556, tmp_pxl_out_557, tmp_pxl_out_558, 
tmp_pxl_out_559, tmp_pxl_out_560, tmp_pxl_out_561, tmp_pxl_out_562, tmp_pxl_out_563, tmp_pxl_out_564, tmp_pxl_out_565, tmp_pxl_out_566, tmp_pxl_out_567, 
tmp_pxl_out_568, tmp_pxl_out_569, tmp_pxl_out_570, tmp_pxl_out_571, tmp_pxl_out_572, tmp_pxl_out_573, tmp_pxl_out_574, tmp_pxl_out_575, tmp_pxl_out_576, 
tmp_pxl_out_577, tmp_pxl_out_578, tmp_pxl_out_579, tmp_pxl_out_580, tmp_pxl_out_581, tmp_pxl_out_582, tmp_pxl_out_583, tmp_pxl_out_584, tmp_pxl_out_585, 
tmp_pxl_out_586, tmp_pxl_out_587, tmp_pxl_out_588, tmp_pxl_out_589, tmp_pxl_out_590, tmp_pxl_out_591, tmp_pxl_out_592, tmp_pxl_out_593, tmp_pxl_out_594, 
tmp_pxl_out_595, tmp_pxl_out_596, tmp_pxl_out_597, tmp_pxl_out_598, tmp_pxl_out_599, tmp_pxl_out_600, tmp_pxl_out_601, tmp_pxl_out_602, tmp_pxl_out_603, 
tmp_pxl_out_604, tmp_pxl_out_605, tmp_pxl_out_606, tmp_pxl_out_607, tmp_pxl_out_608, tmp_pxl_out_609, tmp_pxl_out_610, tmp_pxl_out_611, tmp_pxl_out_612, 
tmp_pxl_out_613, tmp_pxl_out_614, tmp_pxl_out_615, tmp_pxl_out_616, tmp_pxl_out_617, tmp_pxl_out_618, tmp_pxl_out_619, tmp_pxl_out_620, tmp_pxl_out_621, 
tmp_pxl_out_622, tmp_pxl_out_623, tmp_pxl_out_624, tmp_pxl_out_625, tmp_pxl_out_626, tmp_pxl_out_627, tmp_pxl_out_628, tmp_pxl_out_629, tmp_pxl_out_630, 
tmp_pxl_out_631, tmp_pxl_out_632, tmp_pxl_out_633, tmp_pxl_out_634, tmp_pxl_out_635, tmp_pxl_out_636, tmp_pxl_out_637, tmp_pxl_out_638, tmp_pxl_out_639, 
tmp_pxl_out_640, tmp_pxl_out_641, tmp_pxl_out_642, tmp_pxl_out_643, tmp_pxl_out_644, tmp_pxl_out_645, tmp_pxl_out_646, tmp_pxl_out_647, tmp_pxl_out_648, 
tmp_pxl_out_649, tmp_pxl_out_650, tmp_pxl_out_651, tmp_pxl_out_652, tmp_pxl_out_653, tmp_pxl_out_654, tmp_pxl_out_655, tmp_pxl_out_656, tmp_pxl_out_657, 
tmp_pxl_out_658, tmp_pxl_out_659, tmp_pxl_out_660, tmp_pxl_out_661, tmp_pxl_out_662, tmp_pxl_out_663, tmp_pxl_out_664, tmp_pxl_out_665, tmp_pxl_out_666, 
tmp_pxl_out_667, tmp_pxl_out_668, tmp_pxl_out_669, tmp_pxl_out_670, tmp_pxl_out_671, tmp_pxl_out_672, tmp_pxl_out_673, tmp_pxl_out_674, tmp_pxl_out_675, 
tmp_pxl_out_676, tmp_pxl_out_677, tmp_pxl_out_678, tmp_pxl_out_679, tmp_pxl_out_680, tmp_pxl_out_681, tmp_pxl_out_682, tmp_pxl_out_683, tmp_pxl_out_684, 
tmp_pxl_out_685, tmp_pxl_out_686, tmp_pxl_out_687, tmp_pxl_out_688, tmp_pxl_out_689, tmp_pxl_out_690, tmp_pxl_out_691, tmp_pxl_out_692, tmp_pxl_out_693, 
tmp_pxl_out_694, tmp_pxl_out_695, tmp_pxl_out_696, tmp_pxl_out_697, tmp_pxl_out_698, tmp_pxl_out_699, tmp_pxl_out_700, tmp_pxl_out_701, tmp_pxl_out_702, 
tmp_pxl_out_703, tmp_pxl_out_704, tmp_pxl_out_705, tmp_pxl_out_706, tmp_pxl_out_707, tmp_pxl_out_708, tmp_pxl_out_709, tmp_pxl_out_710, tmp_pxl_out_711, 
tmp_pxl_out_712, tmp_pxl_out_713, tmp_pxl_out_714, tmp_pxl_out_715, tmp_pxl_out_716, tmp_pxl_out_717, tmp_pxl_out_718, tmp_pxl_out_719, tmp_pxl_out_720, 
tmp_pxl_out_721, tmp_pxl_out_722, tmp_pxl_out_723, tmp_pxl_out_724, tmp_pxl_out_725, tmp_pxl_out_726, tmp_pxl_out_727, tmp_pxl_out_728, tmp_pxl_out_729, 
tmp_pxl_out_730, tmp_pxl_out_731, tmp_pxl_out_732, tmp_pxl_out_733, tmp_pxl_out_734, tmp_pxl_out_735, tmp_pxl_out_736, tmp_pxl_out_737, tmp_pxl_out_738, 
tmp_pxl_out_739, tmp_pxl_out_740, tmp_pxl_out_741, tmp_pxl_out_742, tmp_pxl_out_743, tmp_pxl_out_744, tmp_pxl_out_745, tmp_pxl_out_746, tmp_pxl_out_747, 
tmp_pxl_out_748, tmp_pxl_out_749, tmp_pxl_out_750, tmp_pxl_out_751, tmp_pxl_out_752, tmp_pxl_out_753, tmp_pxl_out_754, tmp_pxl_out_755, tmp_pxl_out_756, 
tmp_pxl_out_757, tmp_pxl_out_758, tmp_pxl_out_759, tmp_pxl_out_760, tmp_pxl_out_761, tmp_pxl_out_762, tmp_pxl_out_763, tmp_pxl_out_764, tmp_pxl_out_765, 
tmp_pxl_out_766, tmp_pxl_out_767, tmp_pxl_out_768, tmp_pxl_out_769, tmp_pxl_out_770, tmp_pxl_out_771, tmp_pxl_out_772, tmp_pxl_out_773, tmp_pxl_out_774, 
tmp_pxl_out_775, tmp_pxl_out_776, tmp_pxl_out_777, tmp_pxl_out_778, tmp_pxl_out_779, tmp_pxl_out_780, tmp_pxl_out_781, tmp_pxl_out_782, tmp_pxl_out_783, 
tmp_pxl_out_784, tmp_pxl_out_785, tmp_pxl_out_786, tmp_pxl_out_787, tmp_pxl_out_788, tmp_pxl_out_789, tmp_pxl_out_790, tmp_pxl_out_791, tmp_pxl_out_792, 
tmp_pxl_out_793, tmp_pxl_out_794, tmp_pxl_out_795, tmp_pxl_out_796, tmp_pxl_out_797, tmp_pxl_out_798, tmp_pxl_out_799, tmp_pxl_out_800, tmp_pxl_out_801, 
tmp_pxl_out_802, tmp_pxl_out_803, tmp_pxl_out_804, tmp_pxl_out_805, tmp_pxl_out_806, tmp_pxl_out_807, tmp_pxl_out_808, tmp_pxl_out_809, tmp_pxl_out_810, 
tmp_pxl_out_811, tmp_pxl_out_812, tmp_pxl_out_813, tmp_pxl_out_814, tmp_pxl_out_815, tmp_pxl_out_816, tmp_pxl_out_817, tmp_pxl_out_818, tmp_pxl_out_819, 
tmp_pxl_out_820, tmp_pxl_out_821, tmp_pxl_out_822, tmp_pxl_out_823, tmp_pxl_out_824, tmp_pxl_out_825, tmp_pxl_out_826, tmp_pxl_out_827, tmp_pxl_out_828, 
tmp_pxl_out_829, tmp_pxl_out_830, tmp_pxl_out_831, tmp_pxl_out_832, tmp_pxl_out_833, tmp_pxl_out_834, tmp_pxl_out_835, tmp_pxl_out_836, tmp_pxl_out_837, 
tmp_pxl_out_838, tmp_pxl_out_839, tmp_pxl_out_840, tmp_pxl_out_841, tmp_pxl_out_842, tmp_pxl_out_843, tmp_pxl_out_844, tmp_pxl_out_845, tmp_pxl_out_846, 
tmp_pxl_out_847, tmp_pxl_out_848, tmp_pxl_out_849, tmp_pxl_out_850, tmp_pxl_out_851, tmp_pxl_out_852, tmp_pxl_out_853, tmp_pxl_out_854, tmp_pxl_out_855, 
tmp_pxl_out_856, tmp_pxl_out_857, tmp_pxl_out_858, tmp_pxl_out_859, tmp_pxl_out_860, tmp_pxl_out_861, tmp_pxl_out_862, tmp_pxl_out_863, tmp_pxl_out_864, 
tmp_pxl_out_865, tmp_pxl_out_866, tmp_pxl_out_867, tmp_pxl_out_868, tmp_pxl_out_869, tmp_pxl_out_870, tmp_pxl_out_871, tmp_pxl_out_872, tmp_pxl_out_873, 
tmp_pxl_out_874, tmp_pxl_out_875, tmp_pxl_out_876, tmp_pxl_out_877, tmp_pxl_out_878, tmp_pxl_out_879, tmp_pxl_out_880, tmp_pxl_out_881, tmp_pxl_out_882, 
tmp_pxl_out_883, tmp_pxl_out_884, tmp_pxl_out_885, tmp_pxl_out_886, tmp_pxl_out_887, tmp_pxl_out_888, tmp_pxl_out_889, tmp_pxl_out_890, tmp_pxl_out_891, 
tmp_pxl_out_892, tmp_pxl_out_893, tmp_pxl_out_894, tmp_pxl_out_895, tmp_pxl_out_896, tmp_pxl_out_897, tmp_pxl_out_898, tmp_pxl_out_899, tmp_pxl_out_900, 
tmp_pxl_out_901, tmp_pxl_out_902, tmp_pxl_out_903, tmp_pxl_out_904, tmp_pxl_out_905, tmp_pxl_out_906, tmp_pxl_out_907, tmp_pxl_out_908, tmp_pxl_out_909, 
tmp_pxl_out_910, tmp_pxl_out_911, tmp_pxl_out_912, tmp_pxl_out_913, tmp_pxl_out_914, tmp_pxl_out_915, tmp_pxl_out_916, tmp_pxl_out_917, tmp_pxl_out_918, 
tmp_pxl_out_919, tmp_pxl_out_920, tmp_pxl_out_921, tmp_pxl_out_922, tmp_pxl_out_923, tmp_pxl_out_924, tmp_pxl_out_925, tmp_pxl_out_926, tmp_pxl_out_927, 
tmp_pxl_out_928, tmp_pxl_out_929, tmp_pxl_out_930, tmp_pxl_out_931, tmp_pxl_out_932, tmp_pxl_out_933, tmp_pxl_out_934, tmp_pxl_out_935, tmp_pxl_out_936, 
tmp_pxl_out_937, tmp_pxl_out_938, tmp_pxl_out_939, tmp_pxl_out_940, tmp_pxl_out_941, tmp_pxl_out_942, tmp_pxl_out_943, tmp_pxl_out_944, tmp_pxl_out_945, 
tmp_pxl_out_946, tmp_pxl_out_947, tmp_pxl_out_948, tmp_pxl_out_949, tmp_pxl_out_950, tmp_pxl_out_951, tmp_pxl_out_952, tmp_pxl_out_953, tmp_pxl_out_954, 
tmp_pxl_out_955, tmp_pxl_out_956, tmp_pxl_out_957, tmp_pxl_out_958, tmp_pxl_out_959, tmp_pxl_out_960, tmp_pxl_out_961, tmp_pxl_out_962, tmp_pxl_out_963, 
tmp_pxl_out_964, tmp_pxl_out_965, tmp_pxl_out_966, tmp_pxl_out_967, tmp_pxl_out_968, tmp_pxl_out_969, tmp_pxl_out_970, tmp_pxl_out_971, tmp_pxl_out_972, 
tmp_pxl_out_973, tmp_pxl_out_974, tmp_pxl_out_975, tmp_pxl_out_976, tmp_pxl_out_977, tmp_pxl_out_978, tmp_pxl_out_979, tmp_pxl_out_980, tmp_pxl_out_981, 
tmp_pxl_out_982, tmp_pxl_out_983, tmp_pxl_out_984, tmp_pxl_out_985, tmp_pxl_out_986, tmp_pxl_out_987, tmp_pxl_out_988, tmp_pxl_out_989, tmp_pxl_out_990, 
tmp_pxl_out_991, tmp_pxl_out_992, tmp_pxl_out_993, tmp_pxl_out_994, tmp_pxl_out_995, tmp_pxl_out_996, tmp_pxl_out_997, tmp_pxl_out_998, tmp_pxl_out_999, 
tmp_pxl_out_1000, tmp_pxl_out_1001, tmp_pxl_out_1002, tmp_pxl_out_1003, tmp_pxl_out_1004, tmp_pxl_out_1005, tmp_pxl_out_1006, tmp_pxl_out_1007, tmp_pxl_out_1008, 
tmp_pxl_out_1009, tmp_pxl_out_1010, tmp_pxl_out_1011, tmp_pxl_out_1012, tmp_pxl_out_1013, tmp_pxl_out_1014, tmp_pxl_out_1015, tmp_pxl_out_1016, tmp_pxl_out_1017, 
tmp_pxl_out_1018, tmp_pxl_out_1019, tmp_pxl_out_1020, tmp_pxl_out_1021, tmp_pxl_out_1022, tmp_pxl_out_1023, tmp_pxl_out_1024, 
                        
tmp_valid_out_1, tmp_valid_out_2, tmp_valid_out_3, tmp_valid_out_4, tmp_valid_out_5, tmp_valid_out_6, tmp_valid_out_7, tmp_valid_out_8, tmp_valid_out_9, 
tmp_valid_out_10, tmp_valid_out_11, tmp_valid_out_12, tmp_valid_out_13, tmp_valid_out_14, tmp_valid_out_15, tmp_valid_out_16, tmp_valid_out_17, tmp_valid_out_18, 
tmp_valid_out_19, tmp_valid_out_20, tmp_valid_out_21, tmp_valid_out_22, tmp_valid_out_23, tmp_valid_out_24, tmp_valid_out_25, tmp_valid_out_26, tmp_valid_out_27, 
tmp_valid_out_28, tmp_valid_out_29, tmp_valid_out_30, tmp_valid_out_31, tmp_valid_out_32, tmp_valid_out_33, tmp_valid_out_34, tmp_valid_out_35, tmp_valid_out_36, 
tmp_valid_out_37, tmp_valid_out_38, tmp_valid_out_39, tmp_valid_out_40, tmp_valid_out_41, tmp_valid_out_42, tmp_valid_out_43, tmp_valid_out_44, tmp_valid_out_45, 
tmp_valid_out_46, tmp_valid_out_47, tmp_valid_out_48, tmp_valid_out_49, tmp_valid_out_50, tmp_valid_out_51, tmp_valid_out_52, tmp_valid_out_53, tmp_valid_out_54, 
tmp_valid_out_55, tmp_valid_out_56, tmp_valid_out_57, tmp_valid_out_58, tmp_valid_out_59, tmp_valid_out_60, tmp_valid_out_61, tmp_valid_out_62, tmp_valid_out_63, 
tmp_valid_out_64, tmp_valid_out_65, tmp_valid_out_66, tmp_valid_out_67, tmp_valid_out_68, tmp_valid_out_69, tmp_valid_out_70, tmp_valid_out_71, tmp_valid_out_72, 
tmp_valid_out_73, tmp_valid_out_74, tmp_valid_out_75, tmp_valid_out_76, tmp_valid_out_77, tmp_valid_out_78, tmp_valid_out_79, tmp_valid_out_80, tmp_valid_out_81, 
tmp_valid_out_82, tmp_valid_out_83, tmp_valid_out_84, tmp_valid_out_85, tmp_valid_out_86, tmp_valid_out_87, tmp_valid_out_88, tmp_valid_out_89, tmp_valid_out_90, 
tmp_valid_out_91, tmp_valid_out_92, tmp_valid_out_93, tmp_valid_out_94, tmp_valid_out_95, tmp_valid_out_96, tmp_valid_out_97, tmp_valid_out_98, tmp_valid_out_99, 
tmp_valid_out_100, tmp_valid_out_101, tmp_valid_out_102, tmp_valid_out_103, tmp_valid_out_104, tmp_valid_out_105, tmp_valid_out_106, tmp_valid_out_107, tmp_valid_out_108, 
tmp_valid_out_109, tmp_valid_out_110, tmp_valid_out_111, tmp_valid_out_112, tmp_valid_out_113, tmp_valid_out_114, tmp_valid_out_115, tmp_valid_out_116, tmp_valid_out_117, 
tmp_valid_out_118, tmp_valid_out_119, tmp_valid_out_120, tmp_valid_out_121, tmp_valid_out_122, tmp_valid_out_123, tmp_valid_out_124, tmp_valid_out_125, tmp_valid_out_126, 
tmp_valid_out_127, tmp_valid_out_128, tmp_valid_out_129, tmp_valid_out_130, tmp_valid_out_131, tmp_valid_out_132, tmp_valid_out_133, tmp_valid_out_134, tmp_valid_out_135, 
tmp_valid_out_136, tmp_valid_out_137, tmp_valid_out_138, tmp_valid_out_139, tmp_valid_out_140, tmp_valid_out_141, tmp_valid_out_142, tmp_valid_out_143, tmp_valid_out_144, 
tmp_valid_out_145, tmp_valid_out_146, tmp_valid_out_147, tmp_valid_out_148, tmp_valid_out_149, tmp_valid_out_150, tmp_valid_out_151, tmp_valid_out_152, tmp_valid_out_153, 
tmp_valid_out_154, tmp_valid_out_155, tmp_valid_out_156, tmp_valid_out_157, tmp_valid_out_158, tmp_valid_out_159, tmp_valid_out_160, tmp_valid_out_161, tmp_valid_out_162, 
tmp_valid_out_163, tmp_valid_out_164, tmp_valid_out_165, tmp_valid_out_166, tmp_valid_out_167, tmp_valid_out_168, tmp_valid_out_169, tmp_valid_out_170, tmp_valid_out_171, 
tmp_valid_out_172, tmp_valid_out_173, tmp_valid_out_174, tmp_valid_out_175, tmp_valid_out_176, tmp_valid_out_177, tmp_valid_out_178, tmp_valid_out_179, tmp_valid_out_180, 
tmp_valid_out_181, tmp_valid_out_182, tmp_valid_out_183, tmp_valid_out_184, tmp_valid_out_185, tmp_valid_out_186, tmp_valid_out_187, tmp_valid_out_188, tmp_valid_out_189, 
tmp_valid_out_190, tmp_valid_out_191, tmp_valid_out_192, tmp_valid_out_193, tmp_valid_out_194, tmp_valid_out_195, tmp_valid_out_196, tmp_valid_out_197, tmp_valid_out_198, 
tmp_valid_out_199, tmp_valid_out_200, tmp_valid_out_201, tmp_valid_out_202, tmp_valid_out_203, tmp_valid_out_204, tmp_valid_out_205, tmp_valid_out_206, tmp_valid_out_207, 
tmp_valid_out_208, tmp_valid_out_209, tmp_valid_out_210, tmp_valid_out_211, tmp_valid_out_212, tmp_valid_out_213, tmp_valid_out_214, tmp_valid_out_215, tmp_valid_out_216, 
tmp_valid_out_217, tmp_valid_out_218, tmp_valid_out_219, tmp_valid_out_220, tmp_valid_out_221, tmp_valid_out_222, tmp_valid_out_223, tmp_valid_out_224, tmp_valid_out_225, 
tmp_valid_out_226, tmp_valid_out_227, tmp_valid_out_228, tmp_valid_out_229, tmp_valid_out_230, tmp_valid_out_231, tmp_valid_out_232, tmp_valid_out_233, tmp_valid_out_234, 
tmp_valid_out_235, tmp_valid_out_236, tmp_valid_out_237, tmp_valid_out_238, tmp_valid_out_239, tmp_valid_out_240, tmp_valid_out_241, tmp_valid_out_242, tmp_valid_out_243, 
tmp_valid_out_244, tmp_valid_out_245, tmp_valid_out_246, tmp_valid_out_247, tmp_valid_out_248, tmp_valid_out_249, tmp_valid_out_250, tmp_valid_out_251, tmp_valid_out_252, 
tmp_valid_out_253, tmp_valid_out_254, tmp_valid_out_255, tmp_valid_out_256, tmp_valid_out_257, tmp_valid_out_258, tmp_valid_out_259, tmp_valid_out_260, tmp_valid_out_261, 
tmp_valid_out_262, tmp_valid_out_263, tmp_valid_out_264, tmp_valid_out_265, tmp_valid_out_266, tmp_valid_out_267, tmp_valid_out_268, tmp_valid_out_269, tmp_valid_out_270, 
tmp_valid_out_271, tmp_valid_out_272, tmp_valid_out_273, tmp_valid_out_274, tmp_valid_out_275, tmp_valid_out_276, tmp_valid_out_277, tmp_valid_out_278, tmp_valid_out_279, 
tmp_valid_out_280, tmp_valid_out_281, tmp_valid_out_282, tmp_valid_out_283, tmp_valid_out_284, tmp_valid_out_285, tmp_valid_out_286, tmp_valid_out_287, tmp_valid_out_288, 
tmp_valid_out_289, tmp_valid_out_290, tmp_valid_out_291, tmp_valid_out_292, tmp_valid_out_293, tmp_valid_out_294, tmp_valid_out_295, tmp_valid_out_296, tmp_valid_out_297, 
tmp_valid_out_298, tmp_valid_out_299, tmp_valid_out_300, tmp_valid_out_301, tmp_valid_out_302, tmp_valid_out_303, tmp_valid_out_304, tmp_valid_out_305, tmp_valid_out_306, 
tmp_valid_out_307, tmp_valid_out_308, tmp_valid_out_309, tmp_valid_out_310, tmp_valid_out_311, tmp_valid_out_312, tmp_valid_out_313, tmp_valid_out_314, tmp_valid_out_315, 
tmp_valid_out_316, tmp_valid_out_317, tmp_valid_out_318, tmp_valid_out_319, tmp_valid_out_320, tmp_valid_out_321, tmp_valid_out_322, tmp_valid_out_323, tmp_valid_out_324, 
tmp_valid_out_325, tmp_valid_out_326, tmp_valid_out_327, tmp_valid_out_328, tmp_valid_out_329, tmp_valid_out_330, tmp_valid_out_331, tmp_valid_out_332, tmp_valid_out_333, 
tmp_valid_out_334, tmp_valid_out_335, tmp_valid_out_336, tmp_valid_out_337, tmp_valid_out_338, tmp_valid_out_339, tmp_valid_out_340, tmp_valid_out_341, tmp_valid_out_342, 
tmp_valid_out_343, tmp_valid_out_344, tmp_valid_out_345, tmp_valid_out_346, tmp_valid_out_347, tmp_valid_out_348, tmp_valid_out_349, tmp_valid_out_350, tmp_valid_out_351, 
tmp_valid_out_352, tmp_valid_out_353, tmp_valid_out_354, tmp_valid_out_355, tmp_valid_out_356, tmp_valid_out_357, tmp_valid_out_358, tmp_valid_out_359, tmp_valid_out_360, 
tmp_valid_out_361, tmp_valid_out_362, tmp_valid_out_363, tmp_valid_out_364, tmp_valid_out_365, tmp_valid_out_366, tmp_valid_out_367, tmp_valid_out_368, tmp_valid_out_369, 
tmp_valid_out_370, tmp_valid_out_371, tmp_valid_out_372, tmp_valid_out_373, tmp_valid_out_374, tmp_valid_out_375, tmp_valid_out_376, tmp_valid_out_377, tmp_valid_out_378, 
tmp_valid_out_379, tmp_valid_out_380, tmp_valid_out_381, tmp_valid_out_382, tmp_valid_out_383, tmp_valid_out_384, tmp_valid_out_385, tmp_valid_out_386, tmp_valid_out_387, 
tmp_valid_out_388, tmp_valid_out_389, tmp_valid_out_390, tmp_valid_out_391, tmp_valid_out_392, tmp_valid_out_393, tmp_valid_out_394, tmp_valid_out_395, tmp_valid_out_396, 
tmp_valid_out_397, tmp_valid_out_398, tmp_valid_out_399, tmp_valid_out_400, tmp_valid_out_401, tmp_valid_out_402, tmp_valid_out_403, tmp_valid_out_404, tmp_valid_out_405, 
tmp_valid_out_406, tmp_valid_out_407, tmp_valid_out_408, tmp_valid_out_409, tmp_valid_out_410, tmp_valid_out_411, tmp_valid_out_412, tmp_valid_out_413, tmp_valid_out_414, 
tmp_valid_out_415, tmp_valid_out_416, tmp_valid_out_417, tmp_valid_out_418, tmp_valid_out_419, tmp_valid_out_420, tmp_valid_out_421, tmp_valid_out_422, tmp_valid_out_423, 
tmp_valid_out_424, tmp_valid_out_425, tmp_valid_out_426, tmp_valid_out_427, tmp_valid_out_428, tmp_valid_out_429, tmp_valid_out_430, tmp_valid_out_431, tmp_valid_out_432, 
tmp_valid_out_433, tmp_valid_out_434, tmp_valid_out_435, tmp_valid_out_436, tmp_valid_out_437, tmp_valid_out_438, tmp_valid_out_439, tmp_valid_out_440, tmp_valid_out_441, 
tmp_valid_out_442, tmp_valid_out_443, tmp_valid_out_444, tmp_valid_out_445, tmp_valid_out_446, tmp_valid_out_447, tmp_valid_out_448, tmp_valid_out_449, tmp_valid_out_450, 
tmp_valid_out_451, tmp_valid_out_452, tmp_valid_out_453, tmp_valid_out_454, tmp_valid_out_455, tmp_valid_out_456, tmp_valid_out_457, tmp_valid_out_458, tmp_valid_out_459, 
tmp_valid_out_460, tmp_valid_out_461, tmp_valid_out_462, tmp_valid_out_463, tmp_valid_out_464, tmp_valid_out_465, tmp_valid_out_466, tmp_valid_out_467, tmp_valid_out_468, 
tmp_valid_out_469, tmp_valid_out_470, tmp_valid_out_471, tmp_valid_out_472, tmp_valid_out_473, tmp_valid_out_474, tmp_valid_out_475, tmp_valid_out_476, tmp_valid_out_477, 
tmp_valid_out_478, tmp_valid_out_479, tmp_valid_out_480, tmp_valid_out_481, tmp_valid_out_482, tmp_valid_out_483, tmp_valid_out_484, tmp_valid_out_485, tmp_valid_out_486, 
tmp_valid_out_487, tmp_valid_out_488, tmp_valid_out_489, tmp_valid_out_490, tmp_valid_out_491, tmp_valid_out_492, tmp_valid_out_493, tmp_valid_out_494, tmp_valid_out_495, 
tmp_valid_out_496, tmp_valid_out_497, tmp_valid_out_498, tmp_valid_out_499, tmp_valid_out_500, tmp_valid_out_501, tmp_valid_out_502, tmp_valid_out_503, tmp_valid_out_504, 
tmp_valid_out_505, tmp_valid_out_506, tmp_valid_out_507, tmp_valid_out_508, tmp_valid_out_509, tmp_valid_out_510, tmp_valid_out_511, tmp_valid_out_512, tmp_valid_out_513, 
tmp_valid_out_514, tmp_valid_out_515, tmp_valid_out_516, tmp_valid_out_517, tmp_valid_out_518, tmp_valid_out_519, tmp_valid_out_520, tmp_valid_out_521, tmp_valid_out_522, 
tmp_valid_out_523, tmp_valid_out_524, tmp_valid_out_525, tmp_valid_out_526, tmp_valid_out_527, tmp_valid_out_528, tmp_valid_out_529, tmp_valid_out_530, tmp_valid_out_531, 
tmp_valid_out_532, tmp_valid_out_533, tmp_valid_out_534, tmp_valid_out_535, tmp_valid_out_536, tmp_valid_out_537, tmp_valid_out_538, tmp_valid_out_539, tmp_valid_out_540, 
tmp_valid_out_541, tmp_valid_out_542, tmp_valid_out_543, tmp_valid_out_544, tmp_valid_out_545, tmp_valid_out_546, tmp_valid_out_547, tmp_valid_out_548, tmp_valid_out_549, 
tmp_valid_out_550, tmp_valid_out_551, tmp_valid_out_552, tmp_valid_out_553, tmp_valid_out_554, tmp_valid_out_555, tmp_valid_out_556, tmp_valid_out_557, tmp_valid_out_558, 
tmp_valid_out_559, tmp_valid_out_560, tmp_valid_out_561, tmp_valid_out_562, tmp_valid_out_563, tmp_valid_out_564, tmp_valid_out_565, tmp_valid_out_566, tmp_valid_out_567, 
tmp_valid_out_568, tmp_valid_out_569, tmp_valid_out_570, tmp_valid_out_571, tmp_valid_out_572, tmp_valid_out_573, tmp_valid_out_574, tmp_valid_out_575, tmp_valid_out_576, 
tmp_valid_out_577, tmp_valid_out_578, tmp_valid_out_579, tmp_valid_out_580, tmp_valid_out_581, tmp_valid_out_582, tmp_valid_out_583, tmp_valid_out_584, tmp_valid_out_585, 
tmp_valid_out_586, tmp_valid_out_587, tmp_valid_out_588, tmp_valid_out_589, tmp_valid_out_590, tmp_valid_out_591, tmp_valid_out_592, tmp_valid_out_593, tmp_valid_out_594, 
tmp_valid_out_595, tmp_valid_out_596, tmp_valid_out_597, tmp_valid_out_598, tmp_valid_out_599, tmp_valid_out_600, tmp_valid_out_601, tmp_valid_out_602, tmp_valid_out_603, 
tmp_valid_out_604, tmp_valid_out_605, tmp_valid_out_606, tmp_valid_out_607, tmp_valid_out_608, tmp_valid_out_609, tmp_valid_out_610, tmp_valid_out_611, tmp_valid_out_612, 
tmp_valid_out_613, tmp_valid_out_614, tmp_valid_out_615, tmp_valid_out_616, tmp_valid_out_617, tmp_valid_out_618, tmp_valid_out_619, tmp_valid_out_620, tmp_valid_out_621, 
tmp_valid_out_622, tmp_valid_out_623, tmp_valid_out_624, tmp_valid_out_625, tmp_valid_out_626, tmp_valid_out_627, tmp_valid_out_628, tmp_valid_out_629, tmp_valid_out_630, 
tmp_valid_out_631, tmp_valid_out_632, tmp_valid_out_633, tmp_valid_out_634, tmp_valid_out_635, tmp_valid_out_636, tmp_valid_out_637, tmp_valid_out_638, tmp_valid_out_639, 
tmp_valid_out_640, tmp_valid_out_641, tmp_valid_out_642, tmp_valid_out_643, tmp_valid_out_644, tmp_valid_out_645, tmp_valid_out_646, tmp_valid_out_647, tmp_valid_out_648, 
tmp_valid_out_649, tmp_valid_out_650, tmp_valid_out_651, tmp_valid_out_652, tmp_valid_out_653, tmp_valid_out_654, tmp_valid_out_655, tmp_valid_out_656, tmp_valid_out_657, 
tmp_valid_out_658, tmp_valid_out_659, tmp_valid_out_660, tmp_valid_out_661, tmp_valid_out_662, tmp_valid_out_663, tmp_valid_out_664, tmp_valid_out_665, tmp_valid_out_666, 
tmp_valid_out_667, tmp_valid_out_668, tmp_valid_out_669, tmp_valid_out_670, tmp_valid_out_671, tmp_valid_out_672, tmp_valid_out_673, tmp_valid_out_674, tmp_valid_out_675, 
tmp_valid_out_676, tmp_valid_out_677, tmp_valid_out_678, tmp_valid_out_679, tmp_valid_out_680, tmp_valid_out_681, tmp_valid_out_682, tmp_valid_out_683, tmp_valid_out_684, 
tmp_valid_out_685, tmp_valid_out_686, tmp_valid_out_687, tmp_valid_out_688, tmp_valid_out_689, tmp_valid_out_690, tmp_valid_out_691, tmp_valid_out_692, tmp_valid_out_693, 
tmp_valid_out_694, tmp_valid_out_695, tmp_valid_out_696, tmp_valid_out_697, tmp_valid_out_698, tmp_valid_out_699, tmp_valid_out_700, tmp_valid_out_701, tmp_valid_out_702, 
tmp_valid_out_703, tmp_valid_out_704, tmp_valid_out_705, tmp_valid_out_706, tmp_valid_out_707, tmp_valid_out_708, tmp_valid_out_709, tmp_valid_out_710, tmp_valid_out_711, 
tmp_valid_out_712, tmp_valid_out_713, tmp_valid_out_714, tmp_valid_out_715, tmp_valid_out_716, tmp_valid_out_717, tmp_valid_out_718, tmp_valid_out_719, tmp_valid_out_720, 
tmp_valid_out_721, tmp_valid_out_722, tmp_valid_out_723, tmp_valid_out_724, tmp_valid_out_725, tmp_valid_out_726, tmp_valid_out_727, tmp_valid_out_728, tmp_valid_out_729, 
tmp_valid_out_730, tmp_valid_out_731, tmp_valid_out_732, tmp_valid_out_733, tmp_valid_out_734, tmp_valid_out_735, tmp_valid_out_736, tmp_valid_out_737, tmp_valid_out_738, 
tmp_valid_out_739, tmp_valid_out_740, tmp_valid_out_741, tmp_valid_out_742, tmp_valid_out_743, tmp_valid_out_744, tmp_valid_out_745, tmp_valid_out_746, tmp_valid_out_747, 
tmp_valid_out_748, tmp_valid_out_749, tmp_valid_out_750, tmp_valid_out_751, tmp_valid_out_752, tmp_valid_out_753, tmp_valid_out_754, tmp_valid_out_755, tmp_valid_out_756, 
tmp_valid_out_757, tmp_valid_out_758, tmp_valid_out_759, tmp_valid_out_760, tmp_valid_out_761, tmp_valid_out_762, tmp_valid_out_763, tmp_valid_out_764, tmp_valid_out_765, 
tmp_valid_out_766, tmp_valid_out_767, tmp_valid_out_768, tmp_valid_out_769, tmp_valid_out_770, tmp_valid_out_771, tmp_valid_out_772, tmp_valid_out_773, tmp_valid_out_774, 
tmp_valid_out_775, tmp_valid_out_776, tmp_valid_out_777, tmp_valid_out_778, tmp_valid_out_779, tmp_valid_out_780, tmp_valid_out_781, tmp_valid_out_782, tmp_valid_out_783, 
tmp_valid_out_784, tmp_valid_out_785, tmp_valid_out_786, tmp_valid_out_787, tmp_valid_out_788, tmp_valid_out_789, tmp_valid_out_790, tmp_valid_out_791, tmp_valid_out_792, 
tmp_valid_out_793, tmp_valid_out_794, tmp_valid_out_795, tmp_valid_out_796, tmp_valid_out_797, tmp_valid_out_798, tmp_valid_out_799, tmp_valid_out_800, tmp_valid_out_801, 
tmp_valid_out_802, tmp_valid_out_803, tmp_valid_out_804, tmp_valid_out_805, tmp_valid_out_806, tmp_valid_out_807, tmp_valid_out_808, tmp_valid_out_809, tmp_valid_out_810, 
tmp_valid_out_811, tmp_valid_out_812, tmp_valid_out_813, tmp_valid_out_814, tmp_valid_out_815, tmp_valid_out_816, tmp_valid_out_817, tmp_valid_out_818, tmp_valid_out_819, 
tmp_valid_out_820, tmp_valid_out_821, tmp_valid_out_822, tmp_valid_out_823, tmp_valid_out_824, tmp_valid_out_825, tmp_valid_out_826, tmp_valid_out_827, tmp_valid_out_828, 
tmp_valid_out_829, tmp_valid_out_830, tmp_valid_out_831, tmp_valid_out_832, tmp_valid_out_833, tmp_valid_out_834, tmp_valid_out_835, tmp_valid_out_836, tmp_valid_out_837, 
tmp_valid_out_838, tmp_valid_out_839, tmp_valid_out_840, tmp_valid_out_841, tmp_valid_out_842, tmp_valid_out_843, tmp_valid_out_844, tmp_valid_out_845, tmp_valid_out_846, 
tmp_valid_out_847, tmp_valid_out_848, tmp_valid_out_849, tmp_valid_out_850, tmp_valid_out_851, tmp_valid_out_852, tmp_valid_out_853, tmp_valid_out_854, tmp_valid_out_855, 
tmp_valid_out_856, tmp_valid_out_857, tmp_valid_out_858, tmp_valid_out_859, tmp_valid_out_860, tmp_valid_out_861, tmp_valid_out_862, tmp_valid_out_863, tmp_valid_out_864, 
tmp_valid_out_865, tmp_valid_out_866, tmp_valid_out_867, tmp_valid_out_868, tmp_valid_out_869, tmp_valid_out_870, tmp_valid_out_871, tmp_valid_out_872, tmp_valid_out_873, 
tmp_valid_out_874, tmp_valid_out_875, tmp_valid_out_876, tmp_valid_out_877, tmp_valid_out_878, tmp_valid_out_879, tmp_valid_out_880, tmp_valid_out_881, tmp_valid_out_882, 
tmp_valid_out_883, tmp_valid_out_884, tmp_valid_out_885, tmp_valid_out_886, tmp_valid_out_887, tmp_valid_out_888, tmp_valid_out_889, tmp_valid_out_890, tmp_valid_out_891, 
tmp_valid_out_892, tmp_valid_out_893, tmp_valid_out_894, tmp_valid_out_895, tmp_valid_out_896, tmp_valid_out_897, tmp_valid_out_898, tmp_valid_out_899, tmp_valid_out_900, 
tmp_valid_out_901, tmp_valid_out_902, tmp_valid_out_903, tmp_valid_out_904, tmp_valid_out_905, tmp_valid_out_906, tmp_valid_out_907, tmp_valid_out_908, tmp_valid_out_909, 
tmp_valid_out_910, tmp_valid_out_911, tmp_valid_out_912, tmp_valid_out_913, tmp_valid_out_914, tmp_valid_out_915, tmp_valid_out_916, tmp_valid_out_917, tmp_valid_out_918, 
tmp_valid_out_919, tmp_valid_out_920, tmp_valid_out_921, tmp_valid_out_922, tmp_valid_out_923, tmp_valid_out_924, tmp_valid_out_925, tmp_valid_out_926, tmp_valid_out_927, 
tmp_valid_out_928, tmp_valid_out_929, tmp_valid_out_930, tmp_valid_out_931, tmp_valid_out_932, tmp_valid_out_933, tmp_valid_out_934, tmp_valid_out_935, tmp_valid_out_936, 
tmp_valid_out_937, tmp_valid_out_938, tmp_valid_out_939, tmp_valid_out_940, tmp_valid_out_941, tmp_valid_out_942, tmp_valid_out_943, tmp_valid_out_944, tmp_valid_out_945, 
tmp_valid_out_946, tmp_valid_out_947, tmp_valid_out_948, tmp_valid_out_949, tmp_valid_out_950, tmp_valid_out_951, tmp_valid_out_952, tmp_valid_out_953, tmp_valid_out_954, 
tmp_valid_out_955, tmp_valid_out_956, tmp_valid_out_957, tmp_valid_out_958, tmp_valid_out_959, tmp_valid_out_960, tmp_valid_out_961, tmp_valid_out_962, tmp_valid_out_963, 
tmp_valid_out_964, tmp_valid_out_965, tmp_valid_out_966, tmp_valid_out_967, tmp_valid_out_968, tmp_valid_out_969, tmp_valid_out_970, tmp_valid_out_971, tmp_valid_out_972, 
tmp_valid_out_973, tmp_valid_out_974, tmp_valid_out_975, tmp_valid_out_976, tmp_valid_out_977, tmp_valid_out_978, tmp_valid_out_979, tmp_valid_out_980, tmp_valid_out_981, 
tmp_valid_out_982, tmp_valid_out_983, tmp_valid_out_984, tmp_valid_out_985, tmp_valid_out_986, tmp_valid_out_987, tmp_valid_out_988, tmp_valid_out_989, tmp_valid_out_990, 
tmp_valid_out_991, tmp_valid_out_992, tmp_valid_out_993, tmp_valid_out_994, tmp_valid_out_995, tmp_valid_out_996, tmp_valid_out_997, tmp_valid_out_998, tmp_valid_out_999, 
tmp_valid_out_1000, tmp_valid_out_1001, tmp_valid_out_1002, tmp_valid_out_1003, tmp_valid_out_1004, tmp_valid_out_1005, tmp_valid_out_1006, tmp_valid_out_1007, tmp_valid_out_1008, 
tmp_valid_out_1009, tmp_valid_out_1010, tmp_valid_out_1011, tmp_valid_out_1012, tmp_valid_out_1013, tmp_valid_out_1014, tmp_valid_out_1015, tmp_valid_out_1016, tmp_valid_out_1017, 
tmp_valid_out_1018, tmp_valid_out_1019, tmp_valid_out_1020, tmp_valid_out_1021, tmp_valid_out_1022, tmp_valid_out_1023, tmp_valid_out_1024

	);
	
add_1024to32 #((D-2),DATA_WIDTH) uut2 (

clk, 
reset,

tmp_valid_out_1, tmp_valid_out_2, tmp_valid_out_3, tmp_valid_out_4, tmp_valid_out_5, tmp_valid_out_6, tmp_valid_out_7, tmp_valid_out_8, tmp_valid_out_9, 
tmp_valid_out_10, tmp_valid_out_11, tmp_valid_out_12, tmp_valid_out_13, tmp_valid_out_14, tmp_valid_out_15, tmp_valid_out_16, tmp_valid_out_17, tmp_valid_out_18, 
tmp_valid_out_19, tmp_valid_out_20, tmp_valid_out_21, tmp_valid_out_22, tmp_valid_out_23, tmp_valid_out_24, tmp_valid_out_25, tmp_valid_out_26, tmp_valid_out_27, 
tmp_valid_out_28, tmp_valid_out_29, tmp_valid_out_30, tmp_valid_out_31, tmp_valid_out_32, tmp_valid_out_33, tmp_valid_out_34, tmp_valid_out_35, tmp_valid_out_36, 
tmp_valid_out_37, tmp_valid_out_38, tmp_valid_out_39, tmp_valid_out_40, tmp_valid_out_41, tmp_valid_out_42, tmp_valid_out_43, tmp_valid_out_44, tmp_valid_out_45, 
tmp_valid_out_46, tmp_valid_out_47, tmp_valid_out_48, tmp_valid_out_49, tmp_valid_out_50, tmp_valid_out_51, tmp_valid_out_52, tmp_valid_out_53, tmp_valid_out_54, 
tmp_valid_out_55, tmp_valid_out_56, tmp_valid_out_57, tmp_valid_out_58, tmp_valid_out_59, tmp_valid_out_60, tmp_valid_out_61, tmp_valid_out_62, tmp_valid_out_63, 
tmp_valid_out_64, tmp_valid_out_65, tmp_valid_out_66, tmp_valid_out_67, tmp_valid_out_68, tmp_valid_out_69, tmp_valid_out_70, tmp_valid_out_71, tmp_valid_out_72, 
tmp_valid_out_73, tmp_valid_out_74, tmp_valid_out_75, tmp_valid_out_76, tmp_valid_out_77, tmp_valid_out_78, tmp_valid_out_79, tmp_valid_out_80, tmp_valid_out_81, 
tmp_valid_out_82, tmp_valid_out_83, tmp_valid_out_84, tmp_valid_out_85, tmp_valid_out_86, tmp_valid_out_87, tmp_valid_out_88, tmp_valid_out_89, tmp_valid_out_90, 
tmp_valid_out_91, tmp_valid_out_92, tmp_valid_out_93, tmp_valid_out_94, tmp_valid_out_95, tmp_valid_out_96, tmp_valid_out_97, tmp_valid_out_98, tmp_valid_out_99, 
tmp_valid_out_100, tmp_valid_out_101, tmp_valid_out_102, tmp_valid_out_103, tmp_valid_out_104, tmp_valid_out_105, tmp_valid_out_106, tmp_valid_out_107, tmp_valid_out_108, 
tmp_valid_out_109, tmp_valid_out_110, tmp_valid_out_111, tmp_valid_out_112, tmp_valid_out_113, tmp_valid_out_114, tmp_valid_out_115, tmp_valid_out_116, tmp_valid_out_117, 
tmp_valid_out_118, tmp_valid_out_119, tmp_valid_out_120, tmp_valid_out_121, tmp_valid_out_122, tmp_valid_out_123, tmp_valid_out_124, tmp_valid_out_125, tmp_valid_out_126, 
tmp_valid_out_127, tmp_valid_out_128, tmp_valid_out_129, tmp_valid_out_130, tmp_valid_out_131, tmp_valid_out_132, tmp_valid_out_133, tmp_valid_out_134, tmp_valid_out_135, 
tmp_valid_out_136, tmp_valid_out_137, tmp_valid_out_138, tmp_valid_out_139, tmp_valid_out_140, tmp_valid_out_141, tmp_valid_out_142, tmp_valid_out_143, tmp_valid_out_144, 
tmp_valid_out_145, tmp_valid_out_146, tmp_valid_out_147, tmp_valid_out_148, tmp_valid_out_149, tmp_valid_out_150, tmp_valid_out_151, tmp_valid_out_152, tmp_valid_out_153, 
tmp_valid_out_154, tmp_valid_out_155, tmp_valid_out_156, tmp_valid_out_157, tmp_valid_out_158, tmp_valid_out_159, tmp_valid_out_160, tmp_valid_out_161, tmp_valid_out_162, 
tmp_valid_out_163, tmp_valid_out_164, tmp_valid_out_165, tmp_valid_out_166, tmp_valid_out_167, tmp_valid_out_168, tmp_valid_out_169, tmp_valid_out_170, tmp_valid_out_171, 
tmp_valid_out_172, tmp_valid_out_173, tmp_valid_out_174, tmp_valid_out_175, tmp_valid_out_176, tmp_valid_out_177, tmp_valid_out_178, tmp_valid_out_179, tmp_valid_out_180, 
tmp_valid_out_181, tmp_valid_out_182, tmp_valid_out_183, tmp_valid_out_184, tmp_valid_out_185, tmp_valid_out_186, tmp_valid_out_187, tmp_valid_out_188, tmp_valid_out_189, 
tmp_valid_out_190, tmp_valid_out_191, tmp_valid_out_192, tmp_valid_out_193, tmp_valid_out_194, tmp_valid_out_195, tmp_valid_out_196, tmp_valid_out_197, tmp_valid_out_198, 
tmp_valid_out_199, tmp_valid_out_200, tmp_valid_out_201, tmp_valid_out_202, tmp_valid_out_203, tmp_valid_out_204, tmp_valid_out_205, tmp_valid_out_206, tmp_valid_out_207, 
tmp_valid_out_208, tmp_valid_out_209, tmp_valid_out_210, tmp_valid_out_211, tmp_valid_out_212, tmp_valid_out_213, tmp_valid_out_214, tmp_valid_out_215, tmp_valid_out_216, 
tmp_valid_out_217, tmp_valid_out_218, tmp_valid_out_219, tmp_valid_out_220, tmp_valid_out_221, tmp_valid_out_222, tmp_valid_out_223, tmp_valid_out_224, tmp_valid_out_225, 
tmp_valid_out_226, tmp_valid_out_227, tmp_valid_out_228, tmp_valid_out_229, tmp_valid_out_230, tmp_valid_out_231, tmp_valid_out_232, tmp_valid_out_233, tmp_valid_out_234, 
tmp_valid_out_235, tmp_valid_out_236, tmp_valid_out_237, tmp_valid_out_238, tmp_valid_out_239, tmp_valid_out_240, tmp_valid_out_241, tmp_valid_out_242, tmp_valid_out_243, 
tmp_valid_out_244, tmp_valid_out_245, tmp_valid_out_246, tmp_valid_out_247, tmp_valid_out_248, tmp_valid_out_249, tmp_valid_out_250, tmp_valid_out_251, tmp_valid_out_252, 
tmp_valid_out_253, tmp_valid_out_254, tmp_valid_out_255, tmp_valid_out_256, tmp_valid_out_257, tmp_valid_out_258, tmp_valid_out_259, tmp_valid_out_260, tmp_valid_out_261, 
tmp_valid_out_262, tmp_valid_out_263, tmp_valid_out_264, tmp_valid_out_265, tmp_valid_out_266, tmp_valid_out_267, tmp_valid_out_268, tmp_valid_out_269, tmp_valid_out_270, 
tmp_valid_out_271, tmp_valid_out_272, tmp_valid_out_273, tmp_valid_out_274, tmp_valid_out_275, tmp_valid_out_276, tmp_valid_out_277, tmp_valid_out_278, tmp_valid_out_279, 
tmp_valid_out_280, tmp_valid_out_281, tmp_valid_out_282, tmp_valid_out_283, tmp_valid_out_284, tmp_valid_out_285, tmp_valid_out_286, tmp_valid_out_287, tmp_valid_out_288, 
tmp_valid_out_289, tmp_valid_out_290, tmp_valid_out_291, tmp_valid_out_292, tmp_valid_out_293, tmp_valid_out_294, tmp_valid_out_295, tmp_valid_out_296, tmp_valid_out_297, 
tmp_valid_out_298, tmp_valid_out_299, tmp_valid_out_300, tmp_valid_out_301, tmp_valid_out_302, tmp_valid_out_303, tmp_valid_out_304, tmp_valid_out_305, tmp_valid_out_306, 
tmp_valid_out_307, tmp_valid_out_308, tmp_valid_out_309, tmp_valid_out_310, tmp_valid_out_311, tmp_valid_out_312, tmp_valid_out_313, tmp_valid_out_314, tmp_valid_out_315, 
tmp_valid_out_316, tmp_valid_out_317, tmp_valid_out_318, tmp_valid_out_319, tmp_valid_out_320, tmp_valid_out_321, tmp_valid_out_322, tmp_valid_out_323, tmp_valid_out_324, 
tmp_valid_out_325, tmp_valid_out_326, tmp_valid_out_327, tmp_valid_out_328, tmp_valid_out_329, tmp_valid_out_330, tmp_valid_out_331, tmp_valid_out_332, tmp_valid_out_333, 
tmp_valid_out_334, tmp_valid_out_335, tmp_valid_out_336, tmp_valid_out_337, tmp_valid_out_338, tmp_valid_out_339, tmp_valid_out_340, tmp_valid_out_341, tmp_valid_out_342, 
tmp_valid_out_343, tmp_valid_out_344, tmp_valid_out_345, tmp_valid_out_346, tmp_valid_out_347, tmp_valid_out_348, tmp_valid_out_349, tmp_valid_out_350, tmp_valid_out_351, 
tmp_valid_out_352, tmp_valid_out_353, tmp_valid_out_354, tmp_valid_out_355, tmp_valid_out_356, tmp_valid_out_357, tmp_valid_out_358, tmp_valid_out_359, tmp_valid_out_360, 
tmp_valid_out_361, tmp_valid_out_362, tmp_valid_out_363, tmp_valid_out_364, tmp_valid_out_365, tmp_valid_out_366, tmp_valid_out_367, tmp_valid_out_368, tmp_valid_out_369, 
tmp_valid_out_370, tmp_valid_out_371, tmp_valid_out_372, tmp_valid_out_373, tmp_valid_out_374, tmp_valid_out_375, tmp_valid_out_376, tmp_valid_out_377, tmp_valid_out_378, 
tmp_valid_out_379, tmp_valid_out_380, tmp_valid_out_381, tmp_valid_out_382, tmp_valid_out_383, tmp_valid_out_384, tmp_valid_out_385, tmp_valid_out_386, tmp_valid_out_387, 
tmp_valid_out_388, tmp_valid_out_389, tmp_valid_out_390, tmp_valid_out_391, tmp_valid_out_392, tmp_valid_out_393, tmp_valid_out_394, tmp_valid_out_395, tmp_valid_out_396, 
tmp_valid_out_397, tmp_valid_out_398, tmp_valid_out_399, tmp_valid_out_400, tmp_valid_out_401, tmp_valid_out_402, tmp_valid_out_403, tmp_valid_out_404, tmp_valid_out_405, 
tmp_valid_out_406, tmp_valid_out_407, tmp_valid_out_408, tmp_valid_out_409, tmp_valid_out_410, tmp_valid_out_411, tmp_valid_out_412, tmp_valid_out_413, tmp_valid_out_414, 
tmp_valid_out_415, tmp_valid_out_416, tmp_valid_out_417, tmp_valid_out_418, tmp_valid_out_419, tmp_valid_out_420, tmp_valid_out_421, tmp_valid_out_422, tmp_valid_out_423, 
tmp_valid_out_424, tmp_valid_out_425, tmp_valid_out_426, tmp_valid_out_427, tmp_valid_out_428, tmp_valid_out_429, tmp_valid_out_430, tmp_valid_out_431, tmp_valid_out_432, 
tmp_valid_out_433, tmp_valid_out_434, tmp_valid_out_435, tmp_valid_out_436, tmp_valid_out_437, tmp_valid_out_438, tmp_valid_out_439, tmp_valid_out_440, tmp_valid_out_441, 
tmp_valid_out_442, tmp_valid_out_443, tmp_valid_out_444, tmp_valid_out_445, tmp_valid_out_446, tmp_valid_out_447, tmp_valid_out_448, tmp_valid_out_449, tmp_valid_out_450, 
tmp_valid_out_451, tmp_valid_out_452, tmp_valid_out_453, tmp_valid_out_454, tmp_valid_out_455, tmp_valid_out_456, tmp_valid_out_457, tmp_valid_out_458, tmp_valid_out_459, 
tmp_valid_out_460, tmp_valid_out_461, tmp_valid_out_462, tmp_valid_out_463, tmp_valid_out_464, tmp_valid_out_465, tmp_valid_out_466, tmp_valid_out_467, tmp_valid_out_468, 
tmp_valid_out_469, tmp_valid_out_470, tmp_valid_out_471, tmp_valid_out_472, tmp_valid_out_473, tmp_valid_out_474, tmp_valid_out_475, tmp_valid_out_476, tmp_valid_out_477, 
tmp_valid_out_478, tmp_valid_out_479, tmp_valid_out_480, tmp_valid_out_481, tmp_valid_out_482, tmp_valid_out_483, tmp_valid_out_484, tmp_valid_out_485, tmp_valid_out_486, 
tmp_valid_out_487, tmp_valid_out_488, tmp_valid_out_489, tmp_valid_out_490, tmp_valid_out_491, tmp_valid_out_492, tmp_valid_out_493, tmp_valid_out_494, tmp_valid_out_495, 
tmp_valid_out_496, tmp_valid_out_497, tmp_valid_out_498, tmp_valid_out_499, tmp_valid_out_500, tmp_valid_out_501, tmp_valid_out_502, tmp_valid_out_503, tmp_valid_out_504, 
tmp_valid_out_505, tmp_valid_out_506, tmp_valid_out_507, tmp_valid_out_508, tmp_valid_out_509, tmp_valid_out_510, tmp_valid_out_511, tmp_valid_out_512, tmp_valid_out_513, 
tmp_valid_out_514, tmp_valid_out_515, tmp_valid_out_516, tmp_valid_out_517, tmp_valid_out_518, tmp_valid_out_519, tmp_valid_out_520, tmp_valid_out_521, tmp_valid_out_522, 
tmp_valid_out_523, tmp_valid_out_524, tmp_valid_out_525, tmp_valid_out_526, tmp_valid_out_527, tmp_valid_out_528, tmp_valid_out_529, tmp_valid_out_530, tmp_valid_out_531, 
tmp_valid_out_532, tmp_valid_out_533, tmp_valid_out_534, tmp_valid_out_535, tmp_valid_out_536, tmp_valid_out_537, tmp_valid_out_538, tmp_valid_out_539, tmp_valid_out_540, 
tmp_valid_out_541, tmp_valid_out_542, tmp_valid_out_543, tmp_valid_out_544, tmp_valid_out_545, tmp_valid_out_546, tmp_valid_out_547, tmp_valid_out_548, tmp_valid_out_549, 
tmp_valid_out_550, tmp_valid_out_551, tmp_valid_out_552, tmp_valid_out_553, tmp_valid_out_554, tmp_valid_out_555, tmp_valid_out_556, tmp_valid_out_557, tmp_valid_out_558, 
tmp_valid_out_559, tmp_valid_out_560, tmp_valid_out_561, tmp_valid_out_562, tmp_valid_out_563, tmp_valid_out_564, tmp_valid_out_565, tmp_valid_out_566, tmp_valid_out_567, 
tmp_valid_out_568, tmp_valid_out_569, tmp_valid_out_570, tmp_valid_out_571, tmp_valid_out_572, tmp_valid_out_573, tmp_valid_out_574, tmp_valid_out_575, tmp_valid_out_576, 
tmp_valid_out_577, tmp_valid_out_578, tmp_valid_out_579, tmp_valid_out_580, tmp_valid_out_581, tmp_valid_out_582, tmp_valid_out_583, tmp_valid_out_584, tmp_valid_out_585, 
tmp_valid_out_586, tmp_valid_out_587, tmp_valid_out_588, tmp_valid_out_589, tmp_valid_out_590, tmp_valid_out_591, tmp_valid_out_592, tmp_valid_out_593, tmp_valid_out_594, 
tmp_valid_out_595, tmp_valid_out_596, tmp_valid_out_597, tmp_valid_out_598, tmp_valid_out_599, tmp_valid_out_600, tmp_valid_out_601, tmp_valid_out_602, tmp_valid_out_603, 
tmp_valid_out_604, tmp_valid_out_605, tmp_valid_out_606, tmp_valid_out_607, tmp_valid_out_608, tmp_valid_out_609, tmp_valid_out_610, tmp_valid_out_611, tmp_valid_out_612, 
tmp_valid_out_613, tmp_valid_out_614, tmp_valid_out_615, tmp_valid_out_616, tmp_valid_out_617, tmp_valid_out_618, tmp_valid_out_619, tmp_valid_out_620, tmp_valid_out_621, 
tmp_valid_out_622, tmp_valid_out_623, tmp_valid_out_624, tmp_valid_out_625, tmp_valid_out_626, tmp_valid_out_627, tmp_valid_out_628, tmp_valid_out_629, tmp_valid_out_630, 
tmp_valid_out_631, tmp_valid_out_632, tmp_valid_out_633, tmp_valid_out_634, tmp_valid_out_635, tmp_valid_out_636, tmp_valid_out_637, tmp_valid_out_638, tmp_valid_out_639, 
tmp_valid_out_640, tmp_valid_out_641, tmp_valid_out_642, tmp_valid_out_643, tmp_valid_out_644, tmp_valid_out_645, tmp_valid_out_646, tmp_valid_out_647, tmp_valid_out_648, 
tmp_valid_out_649, tmp_valid_out_650, tmp_valid_out_651, tmp_valid_out_652, tmp_valid_out_653, tmp_valid_out_654, tmp_valid_out_655, tmp_valid_out_656, tmp_valid_out_657, 
tmp_valid_out_658, tmp_valid_out_659, tmp_valid_out_660, tmp_valid_out_661, tmp_valid_out_662, tmp_valid_out_663, tmp_valid_out_664, tmp_valid_out_665, tmp_valid_out_666, 
tmp_valid_out_667, tmp_valid_out_668, tmp_valid_out_669, tmp_valid_out_670, tmp_valid_out_671, tmp_valid_out_672, tmp_valid_out_673, tmp_valid_out_674, tmp_valid_out_675, 
tmp_valid_out_676, tmp_valid_out_677, tmp_valid_out_678, tmp_valid_out_679, tmp_valid_out_680, tmp_valid_out_681, tmp_valid_out_682, tmp_valid_out_683, tmp_valid_out_684, 
tmp_valid_out_685, tmp_valid_out_686, tmp_valid_out_687, tmp_valid_out_688, tmp_valid_out_689, tmp_valid_out_690, tmp_valid_out_691, tmp_valid_out_692, tmp_valid_out_693, 
tmp_valid_out_694, tmp_valid_out_695, tmp_valid_out_696, tmp_valid_out_697, tmp_valid_out_698, tmp_valid_out_699, tmp_valid_out_700, tmp_valid_out_701, tmp_valid_out_702, 
tmp_valid_out_703, tmp_valid_out_704, tmp_valid_out_705, tmp_valid_out_706, tmp_valid_out_707, tmp_valid_out_708, tmp_valid_out_709, tmp_valid_out_710, tmp_valid_out_711, 
tmp_valid_out_712, tmp_valid_out_713, tmp_valid_out_714, tmp_valid_out_715, tmp_valid_out_716, tmp_valid_out_717, tmp_valid_out_718, tmp_valid_out_719, tmp_valid_out_720, 
tmp_valid_out_721, tmp_valid_out_722, tmp_valid_out_723, tmp_valid_out_724, tmp_valid_out_725, tmp_valid_out_726, tmp_valid_out_727, tmp_valid_out_728, tmp_valid_out_729, 
tmp_valid_out_730, tmp_valid_out_731, tmp_valid_out_732, tmp_valid_out_733, tmp_valid_out_734, tmp_valid_out_735, tmp_valid_out_736, tmp_valid_out_737, tmp_valid_out_738, 
tmp_valid_out_739, tmp_valid_out_740, tmp_valid_out_741, tmp_valid_out_742, tmp_valid_out_743, tmp_valid_out_744, tmp_valid_out_745, tmp_valid_out_746, tmp_valid_out_747, 
tmp_valid_out_748, tmp_valid_out_749, tmp_valid_out_750, tmp_valid_out_751, tmp_valid_out_752, tmp_valid_out_753, tmp_valid_out_754, tmp_valid_out_755, tmp_valid_out_756, 
tmp_valid_out_757, tmp_valid_out_758, tmp_valid_out_759, tmp_valid_out_760, tmp_valid_out_761, tmp_valid_out_762, tmp_valid_out_763, tmp_valid_out_764, tmp_valid_out_765, 
tmp_valid_out_766, tmp_valid_out_767, tmp_valid_out_768, tmp_valid_out_769, tmp_valid_out_770, tmp_valid_out_771, tmp_valid_out_772, tmp_valid_out_773, tmp_valid_out_774, 
tmp_valid_out_775, tmp_valid_out_776, tmp_valid_out_777, tmp_valid_out_778, tmp_valid_out_779, tmp_valid_out_780, tmp_valid_out_781, tmp_valid_out_782, tmp_valid_out_783, 
tmp_valid_out_784, tmp_valid_out_785, tmp_valid_out_786, tmp_valid_out_787, tmp_valid_out_788, tmp_valid_out_789, tmp_valid_out_790, tmp_valid_out_791, tmp_valid_out_792, 
tmp_valid_out_793, tmp_valid_out_794, tmp_valid_out_795, tmp_valid_out_796, tmp_valid_out_797, tmp_valid_out_798, tmp_valid_out_799, tmp_valid_out_800, tmp_valid_out_801, 
tmp_valid_out_802, tmp_valid_out_803, tmp_valid_out_804, tmp_valid_out_805, tmp_valid_out_806, tmp_valid_out_807, tmp_valid_out_808, tmp_valid_out_809, tmp_valid_out_810, 
tmp_valid_out_811, tmp_valid_out_812, tmp_valid_out_813, tmp_valid_out_814, tmp_valid_out_815, tmp_valid_out_816, tmp_valid_out_817, tmp_valid_out_818, tmp_valid_out_819, 
tmp_valid_out_820, tmp_valid_out_821, tmp_valid_out_822, tmp_valid_out_823, tmp_valid_out_824, tmp_valid_out_825, tmp_valid_out_826, tmp_valid_out_827, tmp_valid_out_828, 
tmp_valid_out_829, tmp_valid_out_830, tmp_valid_out_831, tmp_valid_out_832, tmp_valid_out_833, tmp_valid_out_834, tmp_valid_out_835, tmp_valid_out_836, tmp_valid_out_837, 
tmp_valid_out_838, tmp_valid_out_839, tmp_valid_out_840, tmp_valid_out_841, tmp_valid_out_842, tmp_valid_out_843, tmp_valid_out_844, tmp_valid_out_845, tmp_valid_out_846, 
tmp_valid_out_847, tmp_valid_out_848, tmp_valid_out_849, tmp_valid_out_850, tmp_valid_out_851, tmp_valid_out_852, tmp_valid_out_853, tmp_valid_out_854, tmp_valid_out_855, 
tmp_valid_out_856, tmp_valid_out_857, tmp_valid_out_858, tmp_valid_out_859, tmp_valid_out_860, tmp_valid_out_861, tmp_valid_out_862, tmp_valid_out_863, tmp_valid_out_864, 
tmp_valid_out_865, tmp_valid_out_866, tmp_valid_out_867, tmp_valid_out_868, tmp_valid_out_869, tmp_valid_out_870, tmp_valid_out_871, tmp_valid_out_872, tmp_valid_out_873, 
tmp_valid_out_874, tmp_valid_out_875, tmp_valid_out_876, tmp_valid_out_877, tmp_valid_out_878, tmp_valid_out_879, tmp_valid_out_880, tmp_valid_out_881, tmp_valid_out_882, 
tmp_valid_out_883, tmp_valid_out_884, tmp_valid_out_885, tmp_valid_out_886, tmp_valid_out_887, tmp_valid_out_888, tmp_valid_out_889, tmp_valid_out_890, tmp_valid_out_891, 
tmp_valid_out_892, tmp_valid_out_893, tmp_valid_out_894, tmp_valid_out_895, tmp_valid_out_896, tmp_valid_out_897, tmp_valid_out_898, tmp_valid_out_899, tmp_valid_out_900, 
tmp_valid_out_901, tmp_valid_out_902, tmp_valid_out_903, tmp_valid_out_904, tmp_valid_out_905, tmp_valid_out_906, tmp_valid_out_907, tmp_valid_out_908, tmp_valid_out_909, 
tmp_valid_out_910, tmp_valid_out_911, tmp_valid_out_912, tmp_valid_out_913, tmp_valid_out_914, tmp_valid_out_915, tmp_valid_out_916, tmp_valid_out_917, tmp_valid_out_918, 
tmp_valid_out_919, tmp_valid_out_920, tmp_valid_out_921, tmp_valid_out_922, tmp_valid_out_923, tmp_valid_out_924, tmp_valid_out_925, tmp_valid_out_926, tmp_valid_out_927, 
tmp_valid_out_928, tmp_valid_out_929, tmp_valid_out_930, tmp_valid_out_931, tmp_valid_out_932, tmp_valid_out_933, tmp_valid_out_934, tmp_valid_out_935, tmp_valid_out_936, 
tmp_valid_out_937, tmp_valid_out_938, tmp_valid_out_939, tmp_valid_out_940, tmp_valid_out_941, tmp_valid_out_942, tmp_valid_out_943, tmp_valid_out_944, tmp_valid_out_945, 
tmp_valid_out_946, tmp_valid_out_947, tmp_valid_out_948, tmp_valid_out_949, tmp_valid_out_950, tmp_valid_out_951, tmp_valid_out_952, tmp_valid_out_953, tmp_valid_out_954, 
tmp_valid_out_955, tmp_valid_out_956, tmp_valid_out_957, tmp_valid_out_958, tmp_valid_out_959, tmp_valid_out_960, tmp_valid_out_961, tmp_valid_out_962, tmp_valid_out_963, 
tmp_valid_out_964, tmp_valid_out_965, tmp_valid_out_966, tmp_valid_out_967, tmp_valid_out_968, tmp_valid_out_969, tmp_valid_out_970, tmp_valid_out_971, tmp_valid_out_972, 
tmp_valid_out_973, tmp_valid_out_974, tmp_valid_out_975, tmp_valid_out_976, tmp_valid_out_977, tmp_valid_out_978, tmp_valid_out_979, tmp_valid_out_980, tmp_valid_out_981, 
tmp_valid_out_982, tmp_valid_out_983, tmp_valid_out_984, tmp_valid_out_985, tmp_valid_out_986, tmp_valid_out_987, tmp_valid_out_988, tmp_valid_out_989, tmp_valid_out_990, 
tmp_valid_out_991, tmp_valid_out_992, tmp_valid_out_993, tmp_valid_out_994, tmp_valid_out_995, tmp_valid_out_996, tmp_valid_out_997, tmp_valid_out_998, tmp_valid_out_999, 
tmp_valid_out_1000, tmp_valid_out_1001, tmp_valid_out_1002, tmp_valid_out_1003, tmp_valid_out_1004, tmp_valid_out_1005, tmp_valid_out_1006, tmp_valid_out_1007, tmp_valid_out_1008, 
tmp_valid_out_1009, tmp_valid_out_1010, tmp_valid_out_1011, tmp_valid_out_1012, tmp_valid_out_1013, tmp_valid_out_1014, tmp_valid_out_1015, tmp_valid_out_1016, tmp_valid_out_1017, 
tmp_valid_out_1018, tmp_valid_out_1019, tmp_valid_out_1020, tmp_valid_out_1021, tmp_valid_out_1022, tmp_valid_out_1023, tmp_valid_out_1024, 

tmp_pxl_out_1, tmp_pxl_out_2, tmp_pxl_out_3, tmp_pxl_out_4, tmp_pxl_out_5, tmp_pxl_out_6, tmp_pxl_out_7, tmp_pxl_out_8, tmp_pxl_out_9, 
tmp_pxl_out_10, tmp_pxl_out_11, tmp_pxl_out_12, tmp_pxl_out_13, tmp_pxl_out_14, tmp_pxl_out_15, tmp_pxl_out_16, tmp_pxl_out_17, tmp_pxl_out_18, 
tmp_pxl_out_19, tmp_pxl_out_20, tmp_pxl_out_21, tmp_pxl_out_22, tmp_pxl_out_23, tmp_pxl_out_24, tmp_pxl_out_25, tmp_pxl_out_26, tmp_pxl_out_27, 
tmp_pxl_out_28, tmp_pxl_out_29, tmp_pxl_out_30, tmp_pxl_out_31, tmp_pxl_out_32, tmp_pxl_out_33, tmp_pxl_out_34, tmp_pxl_out_35, tmp_pxl_out_36, 
tmp_pxl_out_37, tmp_pxl_out_38, tmp_pxl_out_39, tmp_pxl_out_40, tmp_pxl_out_41, tmp_pxl_out_42, tmp_pxl_out_43, tmp_pxl_out_44, tmp_pxl_out_45, 
tmp_pxl_out_46, tmp_pxl_out_47, tmp_pxl_out_48, tmp_pxl_out_49, tmp_pxl_out_50, tmp_pxl_out_51, tmp_pxl_out_52, tmp_pxl_out_53, tmp_pxl_out_54, 
tmp_pxl_out_55, tmp_pxl_out_56, tmp_pxl_out_57, tmp_pxl_out_58, tmp_pxl_out_59, tmp_pxl_out_60, tmp_pxl_out_61, tmp_pxl_out_62, tmp_pxl_out_63, 
tmp_pxl_out_64, tmp_pxl_out_65, tmp_pxl_out_66, tmp_pxl_out_67, tmp_pxl_out_68, tmp_pxl_out_69, tmp_pxl_out_70, tmp_pxl_out_71, tmp_pxl_out_72, 
tmp_pxl_out_73, tmp_pxl_out_74, tmp_pxl_out_75, tmp_pxl_out_76, tmp_pxl_out_77, tmp_pxl_out_78, tmp_pxl_out_79, tmp_pxl_out_80, tmp_pxl_out_81, 
tmp_pxl_out_82, tmp_pxl_out_83, tmp_pxl_out_84, tmp_pxl_out_85, tmp_pxl_out_86, tmp_pxl_out_87, tmp_pxl_out_88, tmp_pxl_out_89, tmp_pxl_out_90, 
tmp_pxl_out_91, tmp_pxl_out_92, tmp_pxl_out_93, tmp_pxl_out_94, tmp_pxl_out_95, tmp_pxl_out_96, tmp_pxl_out_97, tmp_pxl_out_98, tmp_pxl_out_99, 
tmp_pxl_out_100, tmp_pxl_out_101, tmp_pxl_out_102, tmp_pxl_out_103, tmp_pxl_out_104, tmp_pxl_out_105, tmp_pxl_out_106, tmp_pxl_out_107, tmp_pxl_out_108, 
tmp_pxl_out_109, tmp_pxl_out_110, tmp_pxl_out_111, tmp_pxl_out_112, tmp_pxl_out_113, tmp_pxl_out_114, tmp_pxl_out_115, tmp_pxl_out_116, tmp_pxl_out_117, 
tmp_pxl_out_118, tmp_pxl_out_119, tmp_pxl_out_120, tmp_pxl_out_121, tmp_pxl_out_122, tmp_pxl_out_123, tmp_pxl_out_124, tmp_pxl_out_125, tmp_pxl_out_126, 
tmp_pxl_out_127, tmp_pxl_out_128, tmp_pxl_out_129, tmp_pxl_out_130, tmp_pxl_out_131, tmp_pxl_out_132, tmp_pxl_out_133, tmp_pxl_out_134, tmp_pxl_out_135, 
tmp_pxl_out_136, tmp_pxl_out_137, tmp_pxl_out_138, tmp_pxl_out_139, tmp_pxl_out_140, tmp_pxl_out_141, tmp_pxl_out_142, tmp_pxl_out_143, tmp_pxl_out_144, 
tmp_pxl_out_145, tmp_pxl_out_146, tmp_pxl_out_147, tmp_pxl_out_148, tmp_pxl_out_149, tmp_pxl_out_150, tmp_pxl_out_151, tmp_pxl_out_152, tmp_pxl_out_153, 
tmp_pxl_out_154, tmp_pxl_out_155, tmp_pxl_out_156, tmp_pxl_out_157, tmp_pxl_out_158, tmp_pxl_out_159, tmp_pxl_out_160, tmp_pxl_out_161, tmp_pxl_out_162, 
tmp_pxl_out_163, tmp_pxl_out_164, tmp_pxl_out_165, tmp_pxl_out_166, tmp_pxl_out_167, tmp_pxl_out_168, tmp_pxl_out_169, tmp_pxl_out_170, tmp_pxl_out_171, 
tmp_pxl_out_172, tmp_pxl_out_173, tmp_pxl_out_174, tmp_pxl_out_175, tmp_pxl_out_176, tmp_pxl_out_177, tmp_pxl_out_178, tmp_pxl_out_179, tmp_pxl_out_180, 
tmp_pxl_out_181, tmp_pxl_out_182, tmp_pxl_out_183, tmp_pxl_out_184, tmp_pxl_out_185, tmp_pxl_out_186, tmp_pxl_out_187, tmp_pxl_out_188, tmp_pxl_out_189, 
tmp_pxl_out_190, tmp_pxl_out_191, tmp_pxl_out_192, tmp_pxl_out_193, tmp_pxl_out_194, tmp_pxl_out_195, tmp_pxl_out_196, tmp_pxl_out_197, tmp_pxl_out_198, 
tmp_pxl_out_199, tmp_pxl_out_200, tmp_pxl_out_201, tmp_pxl_out_202, tmp_pxl_out_203, tmp_pxl_out_204, tmp_pxl_out_205, tmp_pxl_out_206, tmp_pxl_out_207, 
tmp_pxl_out_208, tmp_pxl_out_209, tmp_pxl_out_210, tmp_pxl_out_211, tmp_pxl_out_212, tmp_pxl_out_213, tmp_pxl_out_214, tmp_pxl_out_215, tmp_pxl_out_216, 
tmp_pxl_out_217, tmp_pxl_out_218, tmp_pxl_out_219, tmp_pxl_out_220, tmp_pxl_out_221, tmp_pxl_out_222, tmp_pxl_out_223, tmp_pxl_out_224, tmp_pxl_out_225, 
tmp_pxl_out_226, tmp_pxl_out_227, tmp_pxl_out_228, tmp_pxl_out_229, tmp_pxl_out_230, tmp_pxl_out_231, tmp_pxl_out_232, tmp_pxl_out_233, tmp_pxl_out_234, 
tmp_pxl_out_235, tmp_pxl_out_236, tmp_pxl_out_237, tmp_pxl_out_238, tmp_pxl_out_239, tmp_pxl_out_240, tmp_pxl_out_241, tmp_pxl_out_242, tmp_pxl_out_243, 
tmp_pxl_out_244, tmp_pxl_out_245, tmp_pxl_out_246, tmp_pxl_out_247, tmp_pxl_out_248, tmp_pxl_out_249, tmp_pxl_out_250, tmp_pxl_out_251, tmp_pxl_out_252, 
tmp_pxl_out_253, tmp_pxl_out_254, tmp_pxl_out_255, tmp_pxl_out_256, tmp_pxl_out_257, tmp_pxl_out_258, tmp_pxl_out_259, tmp_pxl_out_260, tmp_pxl_out_261, 
tmp_pxl_out_262, tmp_pxl_out_263, tmp_pxl_out_264, tmp_pxl_out_265, tmp_pxl_out_266, tmp_pxl_out_267, tmp_pxl_out_268, tmp_pxl_out_269, tmp_pxl_out_270, 
tmp_pxl_out_271, tmp_pxl_out_272, tmp_pxl_out_273, tmp_pxl_out_274, tmp_pxl_out_275, tmp_pxl_out_276, tmp_pxl_out_277, tmp_pxl_out_278, tmp_pxl_out_279, 
tmp_pxl_out_280, tmp_pxl_out_281, tmp_pxl_out_282, tmp_pxl_out_283, tmp_pxl_out_284, tmp_pxl_out_285, tmp_pxl_out_286, tmp_pxl_out_287, tmp_pxl_out_288, 
tmp_pxl_out_289, tmp_pxl_out_290, tmp_pxl_out_291, tmp_pxl_out_292, tmp_pxl_out_293, tmp_pxl_out_294, tmp_pxl_out_295, tmp_pxl_out_296, tmp_pxl_out_297, 
tmp_pxl_out_298, tmp_pxl_out_299, tmp_pxl_out_300, tmp_pxl_out_301, tmp_pxl_out_302, tmp_pxl_out_303, tmp_pxl_out_304, tmp_pxl_out_305, tmp_pxl_out_306, 
tmp_pxl_out_307, tmp_pxl_out_308, tmp_pxl_out_309, tmp_pxl_out_310, tmp_pxl_out_311, tmp_pxl_out_312, tmp_pxl_out_313, tmp_pxl_out_314, tmp_pxl_out_315, 
tmp_pxl_out_316, tmp_pxl_out_317, tmp_pxl_out_318, tmp_pxl_out_319, tmp_pxl_out_320, tmp_pxl_out_321, tmp_pxl_out_322, tmp_pxl_out_323, tmp_pxl_out_324, 
tmp_pxl_out_325, tmp_pxl_out_326, tmp_pxl_out_327, tmp_pxl_out_328, tmp_pxl_out_329, tmp_pxl_out_330, tmp_pxl_out_331, tmp_pxl_out_332, tmp_pxl_out_333, 
tmp_pxl_out_334, tmp_pxl_out_335, tmp_pxl_out_336, tmp_pxl_out_337, tmp_pxl_out_338, tmp_pxl_out_339, tmp_pxl_out_340, tmp_pxl_out_341, tmp_pxl_out_342, 
tmp_pxl_out_343, tmp_pxl_out_344, tmp_pxl_out_345, tmp_pxl_out_346, tmp_pxl_out_347, tmp_pxl_out_348, tmp_pxl_out_349, tmp_pxl_out_350, tmp_pxl_out_351, 
tmp_pxl_out_352, tmp_pxl_out_353, tmp_pxl_out_354, tmp_pxl_out_355, tmp_pxl_out_356, tmp_pxl_out_357, tmp_pxl_out_358, tmp_pxl_out_359, tmp_pxl_out_360, 
tmp_pxl_out_361, tmp_pxl_out_362, tmp_pxl_out_363, tmp_pxl_out_364, tmp_pxl_out_365, tmp_pxl_out_366, tmp_pxl_out_367, tmp_pxl_out_368, tmp_pxl_out_369, 
tmp_pxl_out_370, tmp_pxl_out_371, tmp_pxl_out_372, tmp_pxl_out_373, tmp_pxl_out_374, tmp_pxl_out_375, tmp_pxl_out_376, tmp_pxl_out_377, tmp_pxl_out_378, 
tmp_pxl_out_379, tmp_pxl_out_380, tmp_pxl_out_381, tmp_pxl_out_382, tmp_pxl_out_383, tmp_pxl_out_384, tmp_pxl_out_385, tmp_pxl_out_386, tmp_pxl_out_387, 
tmp_pxl_out_388, tmp_pxl_out_389, tmp_pxl_out_390, tmp_pxl_out_391, tmp_pxl_out_392, tmp_pxl_out_393, tmp_pxl_out_394, tmp_pxl_out_395, tmp_pxl_out_396, 
tmp_pxl_out_397, tmp_pxl_out_398, tmp_pxl_out_399, tmp_pxl_out_400, tmp_pxl_out_401, tmp_pxl_out_402, tmp_pxl_out_403, tmp_pxl_out_404, tmp_pxl_out_405, 
tmp_pxl_out_406, tmp_pxl_out_407, tmp_pxl_out_408, tmp_pxl_out_409, tmp_pxl_out_410, tmp_pxl_out_411, tmp_pxl_out_412, tmp_pxl_out_413, tmp_pxl_out_414, 
tmp_pxl_out_415, tmp_pxl_out_416, tmp_pxl_out_417, tmp_pxl_out_418, tmp_pxl_out_419, tmp_pxl_out_420, tmp_pxl_out_421, tmp_pxl_out_422, tmp_pxl_out_423, 
tmp_pxl_out_424, tmp_pxl_out_425, tmp_pxl_out_426, tmp_pxl_out_427, tmp_pxl_out_428, tmp_pxl_out_429, tmp_pxl_out_430, tmp_pxl_out_431, tmp_pxl_out_432, 
tmp_pxl_out_433, tmp_pxl_out_434, tmp_pxl_out_435, tmp_pxl_out_436, tmp_pxl_out_437, tmp_pxl_out_438, tmp_pxl_out_439, tmp_pxl_out_440, tmp_pxl_out_441, 
tmp_pxl_out_442, tmp_pxl_out_443, tmp_pxl_out_444, tmp_pxl_out_445, tmp_pxl_out_446, tmp_pxl_out_447, tmp_pxl_out_448, tmp_pxl_out_449, tmp_pxl_out_450, 
tmp_pxl_out_451, tmp_pxl_out_452, tmp_pxl_out_453, tmp_pxl_out_454, tmp_pxl_out_455, tmp_pxl_out_456, tmp_pxl_out_457, tmp_pxl_out_458, tmp_pxl_out_459, 
tmp_pxl_out_460, tmp_pxl_out_461, tmp_pxl_out_462, tmp_pxl_out_463, tmp_pxl_out_464, tmp_pxl_out_465, tmp_pxl_out_466, tmp_pxl_out_467, tmp_pxl_out_468, 
tmp_pxl_out_469, tmp_pxl_out_470, tmp_pxl_out_471, tmp_pxl_out_472, tmp_pxl_out_473, tmp_pxl_out_474, tmp_pxl_out_475, tmp_pxl_out_476, tmp_pxl_out_477, 
tmp_pxl_out_478, tmp_pxl_out_479, tmp_pxl_out_480, tmp_pxl_out_481, tmp_pxl_out_482, tmp_pxl_out_483, tmp_pxl_out_484, tmp_pxl_out_485, tmp_pxl_out_486, 
tmp_pxl_out_487, tmp_pxl_out_488, tmp_pxl_out_489, tmp_pxl_out_490, tmp_pxl_out_491, tmp_pxl_out_492, tmp_pxl_out_493, tmp_pxl_out_494, tmp_pxl_out_495, 
tmp_pxl_out_496, tmp_pxl_out_497, tmp_pxl_out_498, tmp_pxl_out_499, tmp_pxl_out_500, tmp_pxl_out_501, tmp_pxl_out_502, tmp_pxl_out_503, tmp_pxl_out_504, 
tmp_pxl_out_505, tmp_pxl_out_506, tmp_pxl_out_507, tmp_pxl_out_508, tmp_pxl_out_509, tmp_pxl_out_510, tmp_pxl_out_511, tmp_pxl_out_512, tmp_pxl_out_513, 
tmp_pxl_out_514, tmp_pxl_out_515, tmp_pxl_out_516, tmp_pxl_out_517, tmp_pxl_out_518, tmp_pxl_out_519, tmp_pxl_out_520, tmp_pxl_out_521, tmp_pxl_out_522, 
tmp_pxl_out_523, tmp_pxl_out_524, tmp_pxl_out_525, tmp_pxl_out_526, tmp_pxl_out_527, tmp_pxl_out_528, tmp_pxl_out_529, tmp_pxl_out_530, tmp_pxl_out_531, 
tmp_pxl_out_532, tmp_pxl_out_533, tmp_pxl_out_534, tmp_pxl_out_535, tmp_pxl_out_536, tmp_pxl_out_537, tmp_pxl_out_538, tmp_pxl_out_539, tmp_pxl_out_540, 
tmp_pxl_out_541, tmp_pxl_out_542, tmp_pxl_out_543, tmp_pxl_out_544, tmp_pxl_out_545, tmp_pxl_out_546, tmp_pxl_out_547, tmp_pxl_out_548, tmp_pxl_out_549, 
tmp_pxl_out_550, tmp_pxl_out_551, tmp_pxl_out_552, tmp_pxl_out_553, tmp_pxl_out_554, tmp_pxl_out_555, tmp_pxl_out_556, tmp_pxl_out_557, tmp_pxl_out_558, 
tmp_pxl_out_559, tmp_pxl_out_560, tmp_pxl_out_561, tmp_pxl_out_562, tmp_pxl_out_563, tmp_pxl_out_564, tmp_pxl_out_565, tmp_pxl_out_566, tmp_pxl_out_567, 
tmp_pxl_out_568, tmp_pxl_out_569, tmp_pxl_out_570, tmp_pxl_out_571, tmp_pxl_out_572, tmp_pxl_out_573, tmp_pxl_out_574, tmp_pxl_out_575, tmp_pxl_out_576, 
tmp_pxl_out_577, tmp_pxl_out_578, tmp_pxl_out_579, tmp_pxl_out_580, tmp_pxl_out_581, tmp_pxl_out_582, tmp_pxl_out_583, tmp_pxl_out_584, tmp_pxl_out_585, 
tmp_pxl_out_586, tmp_pxl_out_587, tmp_pxl_out_588, tmp_pxl_out_589, tmp_pxl_out_590, tmp_pxl_out_591, tmp_pxl_out_592, tmp_pxl_out_593, tmp_pxl_out_594, 
tmp_pxl_out_595, tmp_pxl_out_596, tmp_pxl_out_597, tmp_pxl_out_598, tmp_pxl_out_599, tmp_pxl_out_600, tmp_pxl_out_601, tmp_pxl_out_602, tmp_pxl_out_603, 
tmp_pxl_out_604, tmp_pxl_out_605, tmp_pxl_out_606, tmp_pxl_out_607, tmp_pxl_out_608, tmp_pxl_out_609, tmp_pxl_out_610, tmp_pxl_out_611, tmp_pxl_out_612, 
tmp_pxl_out_613, tmp_pxl_out_614, tmp_pxl_out_615, tmp_pxl_out_616, tmp_pxl_out_617, tmp_pxl_out_618, tmp_pxl_out_619, tmp_pxl_out_620, tmp_pxl_out_621, 
tmp_pxl_out_622, tmp_pxl_out_623, tmp_pxl_out_624, tmp_pxl_out_625, tmp_pxl_out_626, tmp_pxl_out_627, tmp_pxl_out_628, tmp_pxl_out_629, tmp_pxl_out_630, 
tmp_pxl_out_631, tmp_pxl_out_632, tmp_pxl_out_633, tmp_pxl_out_634, tmp_pxl_out_635, tmp_pxl_out_636, tmp_pxl_out_637, tmp_pxl_out_638, tmp_pxl_out_639, 
tmp_pxl_out_640, tmp_pxl_out_641, tmp_pxl_out_642, tmp_pxl_out_643, tmp_pxl_out_644, tmp_pxl_out_645, tmp_pxl_out_646, tmp_pxl_out_647, tmp_pxl_out_648, 
tmp_pxl_out_649, tmp_pxl_out_650, tmp_pxl_out_651, tmp_pxl_out_652, tmp_pxl_out_653, tmp_pxl_out_654, tmp_pxl_out_655, tmp_pxl_out_656, tmp_pxl_out_657, 
tmp_pxl_out_658, tmp_pxl_out_659, tmp_pxl_out_660, tmp_pxl_out_661, tmp_pxl_out_662, tmp_pxl_out_663, tmp_pxl_out_664, tmp_pxl_out_665, tmp_pxl_out_666, 
tmp_pxl_out_667, tmp_pxl_out_668, tmp_pxl_out_669, tmp_pxl_out_670, tmp_pxl_out_671, tmp_pxl_out_672, tmp_pxl_out_673, tmp_pxl_out_674, tmp_pxl_out_675, 
tmp_pxl_out_676, tmp_pxl_out_677, tmp_pxl_out_678, tmp_pxl_out_679, tmp_pxl_out_680, tmp_pxl_out_681, tmp_pxl_out_682, tmp_pxl_out_683, tmp_pxl_out_684, 
tmp_pxl_out_685, tmp_pxl_out_686, tmp_pxl_out_687, tmp_pxl_out_688, tmp_pxl_out_689, tmp_pxl_out_690, tmp_pxl_out_691, tmp_pxl_out_692, tmp_pxl_out_693, 
tmp_pxl_out_694, tmp_pxl_out_695, tmp_pxl_out_696, tmp_pxl_out_697, tmp_pxl_out_698, tmp_pxl_out_699, tmp_pxl_out_700, tmp_pxl_out_701, tmp_pxl_out_702, 
tmp_pxl_out_703, tmp_pxl_out_704, tmp_pxl_out_705, tmp_pxl_out_706, tmp_pxl_out_707, tmp_pxl_out_708, tmp_pxl_out_709, tmp_pxl_out_710, tmp_pxl_out_711, 
tmp_pxl_out_712, tmp_pxl_out_713, tmp_pxl_out_714, tmp_pxl_out_715, tmp_pxl_out_716, tmp_pxl_out_717, tmp_pxl_out_718, tmp_pxl_out_719, tmp_pxl_out_720, 
tmp_pxl_out_721, tmp_pxl_out_722, tmp_pxl_out_723, tmp_pxl_out_724, tmp_pxl_out_725, tmp_pxl_out_726, tmp_pxl_out_727, tmp_pxl_out_728, tmp_pxl_out_729, 
tmp_pxl_out_730, tmp_pxl_out_731, tmp_pxl_out_732, tmp_pxl_out_733, tmp_pxl_out_734, tmp_pxl_out_735, tmp_pxl_out_736, tmp_pxl_out_737, tmp_pxl_out_738, 
tmp_pxl_out_739, tmp_pxl_out_740, tmp_pxl_out_741, tmp_pxl_out_742, tmp_pxl_out_743, tmp_pxl_out_744, tmp_pxl_out_745, tmp_pxl_out_746, tmp_pxl_out_747, 
tmp_pxl_out_748, tmp_pxl_out_749, tmp_pxl_out_750, tmp_pxl_out_751, tmp_pxl_out_752, tmp_pxl_out_753, tmp_pxl_out_754, tmp_pxl_out_755, tmp_pxl_out_756, 
tmp_pxl_out_757, tmp_pxl_out_758, tmp_pxl_out_759, tmp_pxl_out_760, tmp_pxl_out_761, tmp_pxl_out_762, tmp_pxl_out_763, tmp_pxl_out_764, tmp_pxl_out_765, 
tmp_pxl_out_766, tmp_pxl_out_767, tmp_pxl_out_768, tmp_pxl_out_769, tmp_pxl_out_770, tmp_pxl_out_771, tmp_pxl_out_772, tmp_pxl_out_773, tmp_pxl_out_774, 
tmp_pxl_out_775, tmp_pxl_out_776, tmp_pxl_out_777, tmp_pxl_out_778, tmp_pxl_out_779, tmp_pxl_out_780, tmp_pxl_out_781, tmp_pxl_out_782, tmp_pxl_out_783, 
tmp_pxl_out_784, tmp_pxl_out_785, tmp_pxl_out_786, tmp_pxl_out_787, tmp_pxl_out_788, tmp_pxl_out_789, tmp_pxl_out_790, tmp_pxl_out_791, tmp_pxl_out_792, 
tmp_pxl_out_793, tmp_pxl_out_794, tmp_pxl_out_795, tmp_pxl_out_796, tmp_pxl_out_797, tmp_pxl_out_798, tmp_pxl_out_799, tmp_pxl_out_800, tmp_pxl_out_801, 
tmp_pxl_out_802, tmp_pxl_out_803, tmp_pxl_out_804, tmp_pxl_out_805, tmp_pxl_out_806, tmp_pxl_out_807, tmp_pxl_out_808, tmp_pxl_out_809, tmp_pxl_out_810, 
tmp_pxl_out_811, tmp_pxl_out_812, tmp_pxl_out_813, tmp_pxl_out_814, tmp_pxl_out_815, tmp_pxl_out_816, tmp_pxl_out_817, tmp_pxl_out_818, tmp_pxl_out_819, 
tmp_pxl_out_820, tmp_pxl_out_821, tmp_pxl_out_822, tmp_pxl_out_823, tmp_pxl_out_824, tmp_pxl_out_825, tmp_pxl_out_826, tmp_pxl_out_827, tmp_pxl_out_828, 
tmp_pxl_out_829, tmp_pxl_out_830, tmp_pxl_out_831, tmp_pxl_out_832, tmp_pxl_out_833, tmp_pxl_out_834, tmp_pxl_out_835, tmp_pxl_out_836, tmp_pxl_out_837, 
tmp_pxl_out_838, tmp_pxl_out_839, tmp_pxl_out_840, tmp_pxl_out_841, tmp_pxl_out_842, tmp_pxl_out_843, tmp_pxl_out_844, tmp_pxl_out_845, tmp_pxl_out_846, 
tmp_pxl_out_847, tmp_pxl_out_848, tmp_pxl_out_849, tmp_pxl_out_850, tmp_pxl_out_851, tmp_pxl_out_852, tmp_pxl_out_853, tmp_pxl_out_854, tmp_pxl_out_855, 
tmp_pxl_out_856, tmp_pxl_out_857, tmp_pxl_out_858, tmp_pxl_out_859, tmp_pxl_out_860, tmp_pxl_out_861, tmp_pxl_out_862, tmp_pxl_out_863, tmp_pxl_out_864, 
tmp_pxl_out_865, tmp_pxl_out_866, tmp_pxl_out_867, tmp_pxl_out_868, tmp_pxl_out_869, tmp_pxl_out_870, tmp_pxl_out_871, tmp_pxl_out_872, tmp_pxl_out_873, 
tmp_pxl_out_874, tmp_pxl_out_875, tmp_pxl_out_876, tmp_pxl_out_877, tmp_pxl_out_878, tmp_pxl_out_879, tmp_pxl_out_880, tmp_pxl_out_881, tmp_pxl_out_882, 
tmp_pxl_out_883, tmp_pxl_out_884, tmp_pxl_out_885, tmp_pxl_out_886, tmp_pxl_out_887, tmp_pxl_out_888, tmp_pxl_out_889, tmp_pxl_out_890, tmp_pxl_out_891, 
tmp_pxl_out_892, tmp_pxl_out_893, tmp_pxl_out_894, tmp_pxl_out_895, tmp_pxl_out_896, tmp_pxl_out_897, tmp_pxl_out_898, tmp_pxl_out_899, tmp_pxl_out_900, 
tmp_pxl_out_901, tmp_pxl_out_902, tmp_pxl_out_903, tmp_pxl_out_904, tmp_pxl_out_905, tmp_pxl_out_906, tmp_pxl_out_907, tmp_pxl_out_908, tmp_pxl_out_909, 
tmp_pxl_out_910, tmp_pxl_out_911, tmp_pxl_out_912, tmp_pxl_out_913, tmp_pxl_out_914, tmp_pxl_out_915, tmp_pxl_out_916, tmp_pxl_out_917, tmp_pxl_out_918, 
tmp_pxl_out_919, tmp_pxl_out_920, tmp_pxl_out_921, tmp_pxl_out_922, tmp_pxl_out_923, tmp_pxl_out_924, tmp_pxl_out_925, tmp_pxl_out_926, tmp_pxl_out_927, 
tmp_pxl_out_928, tmp_pxl_out_929, tmp_pxl_out_930, tmp_pxl_out_931, tmp_pxl_out_932, tmp_pxl_out_933, tmp_pxl_out_934, tmp_pxl_out_935, tmp_pxl_out_936, 
tmp_pxl_out_937, tmp_pxl_out_938, tmp_pxl_out_939, tmp_pxl_out_940, tmp_pxl_out_941, tmp_pxl_out_942, tmp_pxl_out_943, tmp_pxl_out_944, tmp_pxl_out_945, 
tmp_pxl_out_946, tmp_pxl_out_947, tmp_pxl_out_948, tmp_pxl_out_949, tmp_pxl_out_950, tmp_pxl_out_951, tmp_pxl_out_952, tmp_pxl_out_953, tmp_pxl_out_954, 
tmp_pxl_out_955, tmp_pxl_out_956, tmp_pxl_out_957, tmp_pxl_out_958, tmp_pxl_out_959, tmp_pxl_out_960, tmp_pxl_out_961, tmp_pxl_out_962, tmp_pxl_out_963, 
tmp_pxl_out_964, tmp_pxl_out_965, tmp_pxl_out_966, tmp_pxl_out_967, tmp_pxl_out_968, tmp_pxl_out_969, tmp_pxl_out_970, tmp_pxl_out_971, tmp_pxl_out_972, 
tmp_pxl_out_973, tmp_pxl_out_974, tmp_pxl_out_975, tmp_pxl_out_976, tmp_pxl_out_977, tmp_pxl_out_978, tmp_pxl_out_979, tmp_pxl_out_980, tmp_pxl_out_981, 
tmp_pxl_out_982, tmp_pxl_out_983, tmp_pxl_out_984, tmp_pxl_out_985, tmp_pxl_out_986, tmp_pxl_out_987, tmp_pxl_out_988, tmp_pxl_out_989, tmp_pxl_out_990, 
tmp_pxl_out_991, tmp_pxl_out_992, tmp_pxl_out_993, tmp_pxl_out_994, tmp_pxl_out_995, tmp_pxl_out_996, tmp_pxl_out_997, tmp_pxl_out_998, tmp_pxl_out_999, 
tmp_pxl_out_1000, tmp_pxl_out_1001, tmp_pxl_out_1002, tmp_pxl_out_1003, tmp_pxl_out_1004, tmp_pxl_out_1005, tmp_pxl_out_1006, tmp_pxl_out_1007, tmp_pxl_out_1008, 
tmp_pxl_out_1009, tmp_pxl_out_1010, tmp_pxl_out_1011, tmp_pxl_out_1012, tmp_pxl_out_1013, tmp_pxl_out_1014, tmp_pxl_out_1015, tmp_pxl_out_1016, tmp_pxl_out_1017, 
tmp_pxl_out_1018, tmp_pxl_out_1019, tmp_pxl_out_1020, tmp_pxl_out_1021, tmp_pxl_out_1022, tmp_pxl_out_1023, tmp_pxl_out_1024, 

    	                   pxl_out_1 , pxl_out_2 , pxl_out_3 , pxl_out_4 , pxl_out_5 , pxl_out_6 , pxl_out_7 , pxl_out_8 , pxl_out_9 , pxl_out_10,
                        pxl_out_11, pxl_out_12, pxl_out_13, pxl_out_14, pxl_out_15, pxl_out_16, pxl_out_17, pxl_out_18, pxl_out_19, pxl_out_20,
	                      pxl_out_21, pxl_out_22, pxl_out_23, pxl_out_24, pxl_out_25, pxl_out_26, pxl_out_27, pxl_out_28, pxl_out_29, pxl_out_30,
                        pxl_out_31, pxl_out_32,
	                                 
	                      valid_out_1 , valid_out_2 , valid_out_3 , valid_out_4 , valid_out_5 , valid_out_6 , valid_out_7 , valid_out_8 , valid_out_9 , valid_out_10,
                        valid_out_11, valid_out_12, valid_out_13, valid_out_14, valid_out_15, valid_out_16, valid_out_17, valid_out_18, valid_out_19, valid_out_20,
	                      valid_out_21, valid_out_22, valid_out_23, valid_out_24, valid_out_25, valid_out_26, valid_out_27, valid_out_28, valid_out_29, valid_out_30,
                        valid_out_31, valid_out_32
);

endmodule