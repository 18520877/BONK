`timescale 1ns / 1ps
// Convolution Kernel 3x3, Stride = 2, Padding = 0.

module tb_Conv2d_2a_3x3_32;
  parameter data_width = 32;
  parameter D = 9;
  parameter T = D*D;
	parameter C = 10;
	parameter I = 20;
	integer i;
	/*integer j;
	integer g;*/
	
	reg clk;
	reg reset;
	     	reg valid_in_1,  valid_in_2,  valid_in_3,  valid_in_4,  valid_in_5,  valid_in_6,
    	       valid_in_7,  valid_in_8,  valid_in_9,  valid_in_10, valid_in_11, valid_in_12,
    	       valid_in_13, valid_in_14, valid_in_15, valid_in_16, valid_in_17, valid_in_18,
    	       valid_in_19, valid_in_20, valid_in_21, valid_in_22, valid_in_23, valid_in_24,
  	         valid_in_25, valid_in_26, valid_in_27, valid_in_28, valid_in_29, valid_in_30,
    	       valid_in_31, valid_in_32;
    	      
    	  reg [data_width-1:0] pxl_in_1,  pxl_in_2,  pxl_in_3,  pxl_in_4,  pxl_in_5,  pxl_in_6,
    	                       pxl_in_7,  pxl_in_8,  pxl_in_9,  pxl_in_10, pxl_in_11, pxl_in_12,
    	                       pxl_in_13, pxl_in_14, pxl_in_15, pxl_in_16, pxl_in_17, pxl_in_18,
    	                       pxl_in_19, pxl_in_20, pxl_in_21, pxl_in_22, pxl_in_23, pxl_in_24,
    	                       pxl_in_25, pxl_in_26, pxl_in_27, pxl_in_28, pxl_in_29, pxl_in_30,
    	                       pxl_in_31, pxl_in_32;

	
	reg [data_width-1:0]In1[T-1:0];
	reg [data_width-1:0]In2[T-1:0];
	reg [data_width-1:0]In3[T-1:0];
	reg [data_width-1:0]In4[T-1:0];
	reg [data_width-1:0]In5[T-1:0];
	reg [data_width-1:0]In6[T-1:0];
	reg [data_width-1:0]In7[T-1:0];
	reg [data_width-1:0]In8[T-1:0];
	reg [data_width-1:0]In9[T-1:0];
	reg [data_width-1:0]In10[T-1:0];
	reg [data_width-1:0]In11[T-1:0];
	reg [data_width-1:0]In12[T-1:0];
	reg [data_width-1:0]In13[T-1:0];
	reg [data_width-1:0]In14[T-1:0];
	reg [data_width-1:0]In15[T-1:0];
	reg [data_width-1:0]In16[T-1:0];
	reg [data_width-1:0]In17[T-1:0];
	reg [data_width-1:0]In18[T-1:0];
	reg [data_width-1:0]In19[T-1:0];
	reg [data_width-1:0]In20[T-1:0];
	reg [data_width-1:0]In21[T-1:0];
	reg [data_width-1:0]In22[T-1:0];
	reg [data_width-1:0]In23[T-1:0];
	reg [data_width-1:0]In24[T-1:0];
	reg [data_width-1:0]In25[T-1:0];
	reg [data_width-1:0]In26[T-1:0];
	reg [data_width-1:0]In27[T-1:0];
	reg [data_width-1:0]In28[T-1:0];
	reg [data_width-1:0]In29[T-1:0];
	reg [data_width-1:0]In30[T-1:0];
	reg [data_width-1:0]In31[T-1:0];
	reg [data_width-1:0]In32[T-1:0];
	


  wire [data_width-1:0] pxl_out_1,pxl_out_2,pxl_out_3,pxl_out_4,pxl_out_5,pxl_out_6,pxl_out_7,pxl_out_8,pxl_out_9,
pxl_out_10,pxl_out_11,pxl_out_12,pxl_out_13,pxl_out_14,pxl_out_15,pxl_out_16,pxl_out_17,pxl_out_18,
pxl_out_19,pxl_out_20,pxl_out_21,pxl_out_22,pxl_out_23,pxl_out_24,pxl_out_25,pxl_out_26,pxl_out_27,
pxl_out_28,pxl_out_29,pxl_out_30,pxl_out_31,pxl_out_32,pxl_out_33,pxl_out_34,pxl_out_35,pxl_out_36,
pxl_out_37,pxl_out_38,pxl_out_39,pxl_out_40,pxl_out_41,pxl_out_42,pxl_out_43,pxl_out_44,pxl_out_45,
pxl_out_46,pxl_out_47,pxl_out_48,pxl_out_49,pxl_out_50,pxl_out_51,pxl_out_52,pxl_out_53,pxl_out_54,
pxl_out_55,pxl_out_56,pxl_out_57,pxl_out_58,pxl_out_59,pxl_out_60,pxl_out_61,pxl_out_62,pxl_out_63,
pxl_out_64,pxl_out_65,pxl_out_66,pxl_out_67,pxl_out_68,pxl_out_69,pxl_out_70,pxl_out_71,pxl_out_72,
pxl_out_73,pxl_out_74,pxl_out_75,pxl_out_76,pxl_out_77,pxl_out_78,pxl_out_79,pxl_out_80,pxl_out_81,
pxl_out_82,pxl_out_83,pxl_out_84,pxl_out_85,pxl_out_86,pxl_out_87,pxl_out_88,pxl_out_89,pxl_out_90,
pxl_out_91,pxl_out_92,pxl_out_93,pxl_out_94,pxl_out_95,pxl_out_96,pxl_out_97,pxl_out_98,pxl_out_99,
pxl_out_100,pxl_out_101,pxl_out_102,pxl_out_103,pxl_out_104,pxl_out_105,pxl_out_106,pxl_out_107,pxl_out_108,
pxl_out_109,pxl_out_110,pxl_out_111,pxl_out_112,pxl_out_113,pxl_out_114,pxl_out_115,pxl_out_116,pxl_out_117,
pxl_out_118,pxl_out_119,pxl_out_120,pxl_out_121,pxl_out_122,pxl_out_123,pxl_out_124,pxl_out_125,pxl_out_126,
pxl_out_127,pxl_out_128,pxl_out_129,pxl_out_130,pxl_out_131,pxl_out_132,pxl_out_133,pxl_out_134,pxl_out_135,
pxl_out_136,pxl_out_137,pxl_out_138,pxl_out_139,pxl_out_140,pxl_out_141,pxl_out_142,pxl_out_143,pxl_out_144,
pxl_out_145,pxl_out_146,pxl_out_147,pxl_out_148,pxl_out_149,pxl_out_150,pxl_out_151,pxl_out_152,pxl_out_153,
pxl_out_154,pxl_out_155,pxl_out_156,pxl_out_157,pxl_out_158,pxl_out_159,pxl_out_160,pxl_out_161,pxl_out_162,
pxl_out_163,pxl_out_164,pxl_out_165,pxl_out_166,pxl_out_167,pxl_out_168,pxl_out_169,pxl_out_170,pxl_out_171,
pxl_out_172,pxl_out_173,pxl_out_174,pxl_out_175,pxl_out_176,pxl_out_177,pxl_out_178,pxl_out_179,pxl_out_180,
pxl_out_181,pxl_out_182,pxl_out_183,pxl_out_184,pxl_out_185,pxl_out_186,pxl_out_187,pxl_out_188,pxl_out_189,
pxl_out_190,pxl_out_191,pxl_out_192,pxl_out_193,pxl_out_194,pxl_out_195,pxl_out_196,pxl_out_197,pxl_out_198,
pxl_out_199,pxl_out_200,pxl_out_201,pxl_out_202,pxl_out_203,pxl_out_204,pxl_out_205,pxl_out_206,pxl_out_207,
pxl_out_208,pxl_out_209,pxl_out_210,pxl_out_211,pxl_out_212,pxl_out_213,pxl_out_214,pxl_out_215,pxl_out_216,
pxl_out_217,pxl_out_218,pxl_out_219,pxl_out_220,pxl_out_221,pxl_out_222,pxl_out_223,pxl_out_224,pxl_out_225,
pxl_out_226,pxl_out_227,pxl_out_228,pxl_out_229,pxl_out_230,pxl_out_231,pxl_out_232,pxl_out_233,pxl_out_234,
pxl_out_235,pxl_out_236,pxl_out_237,pxl_out_238,pxl_out_239,pxl_out_240,pxl_out_241,pxl_out_242,pxl_out_243,
pxl_out_244,pxl_out_245,pxl_out_246,pxl_out_247,pxl_out_248,pxl_out_249,pxl_out_250,pxl_out_251,pxl_out_252,
pxl_out_253,pxl_out_254,pxl_out_255,pxl_out_256,pxl_out_257,pxl_out_258,pxl_out_259,pxl_out_260,pxl_out_261,
pxl_out_262,pxl_out_263,pxl_out_264,pxl_out_265,pxl_out_266,pxl_out_267,pxl_out_268,pxl_out_269,pxl_out_270,
pxl_out_271,pxl_out_272,pxl_out_273,pxl_out_274,pxl_out_275,pxl_out_276,pxl_out_277,pxl_out_278,pxl_out_279,
pxl_out_280,pxl_out_281,pxl_out_282,pxl_out_283,pxl_out_284,pxl_out_285,pxl_out_286,pxl_out_287,pxl_out_288,
pxl_out_289,pxl_out_290,pxl_out_291,pxl_out_292,pxl_out_293,pxl_out_294,pxl_out_295,pxl_out_296,pxl_out_297,
pxl_out_298,pxl_out_299,pxl_out_300,pxl_out_301,pxl_out_302,pxl_out_303,pxl_out_304,pxl_out_305,pxl_out_306,
pxl_out_307,pxl_out_308,pxl_out_309,pxl_out_310,pxl_out_311,pxl_out_312,pxl_out_313,pxl_out_314,pxl_out_315,
pxl_out_316,pxl_out_317,pxl_out_318,pxl_out_319,pxl_out_320,pxl_out_321,pxl_out_322,pxl_out_323,pxl_out_324,
pxl_out_325,pxl_out_326,pxl_out_327,pxl_out_328,pxl_out_329,pxl_out_330,pxl_out_331,pxl_out_332,pxl_out_333,
pxl_out_334,pxl_out_335,pxl_out_336,pxl_out_337,pxl_out_338,pxl_out_339,pxl_out_340,pxl_out_341,pxl_out_342,
pxl_out_343,pxl_out_344,pxl_out_345,pxl_out_346,pxl_out_347,pxl_out_348,pxl_out_349,pxl_out_350,pxl_out_351,
pxl_out_352,pxl_out_353,pxl_out_354,pxl_out_355,pxl_out_356,pxl_out_357,pxl_out_358,pxl_out_359,pxl_out_360,
pxl_out_361,pxl_out_362,pxl_out_363,pxl_out_364,pxl_out_365,pxl_out_366,pxl_out_367,pxl_out_368,pxl_out_369,
pxl_out_370,pxl_out_371,pxl_out_372,pxl_out_373,pxl_out_374,pxl_out_375,pxl_out_376,pxl_out_377,pxl_out_378,
pxl_out_379,pxl_out_380,pxl_out_381,pxl_out_382,pxl_out_383,pxl_out_384,pxl_out_385,pxl_out_386,pxl_out_387,
pxl_out_388,pxl_out_389,pxl_out_390,pxl_out_391,pxl_out_392,pxl_out_393,pxl_out_394,pxl_out_395,pxl_out_396,
pxl_out_397,pxl_out_398,pxl_out_399,pxl_out_400,pxl_out_401,pxl_out_402,pxl_out_403,pxl_out_404,pxl_out_405,
pxl_out_406,pxl_out_407,pxl_out_408,pxl_out_409,pxl_out_410,pxl_out_411,pxl_out_412,pxl_out_413,pxl_out_414,
pxl_out_415,pxl_out_416,pxl_out_417,pxl_out_418,pxl_out_419,pxl_out_420,pxl_out_421,pxl_out_422,pxl_out_423,
pxl_out_424,pxl_out_425,pxl_out_426,pxl_out_427,pxl_out_428,pxl_out_429,pxl_out_430,pxl_out_431,pxl_out_432,
pxl_out_433,pxl_out_434,pxl_out_435,pxl_out_436,pxl_out_437,pxl_out_438,pxl_out_439,pxl_out_440,pxl_out_441,
pxl_out_442,pxl_out_443,pxl_out_444,pxl_out_445,pxl_out_446,pxl_out_447,pxl_out_448,pxl_out_449,pxl_out_450,
pxl_out_451,pxl_out_452,pxl_out_453,pxl_out_454,pxl_out_455,pxl_out_456,pxl_out_457,pxl_out_458,pxl_out_459,
pxl_out_460,pxl_out_461,pxl_out_462,pxl_out_463,pxl_out_464,pxl_out_465,pxl_out_466,pxl_out_467,pxl_out_468,
pxl_out_469,pxl_out_470,pxl_out_471,pxl_out_472,pxl_out_473,pxl_out_474,pxl_out_475,pxl_out_476,pxl_out_477,
pxl_out_478,pxl_out_479,pxl_out_480,pxl_out_481,pxl_out_482,pxl_out_483,pxl_out_484,pxl_out_485,pxl_out_486,
pxl_out_487,pxl_out_488,pxl_out_489,pxl_out_490,pxl_out_491,pxl_out_492,pxl_out_493,pxl_out_494,pxl_out_495,
pxl_out_496,pxl_out_497,pxl_out_498,pxl_out_499,pxl_out_500,pxl_out_501,pxl_out_502,pxl_out_503,pxl_out_504,
pxl_out_505,pxl_out_506,pxl_out_507,pxl_out_508,pxl_out_509,pxl_out_510,pxl_out_511,pxl_out_512,pxl_out_513,
pxl_out_514,pxl_out_515,pxl_out_516,pxl_out_517,pxl_out_518,pxl_out_519,pxl_out_520,pxl_out_521,pxl_out_522,
pxl_out_523,pxl_out_524,pxl_out_525,pxl_out_526,pxl_out_527,pxl_out_528,pxl_out_529,pxl_out_530,pxl_out_531,
pxl_out_532,pxl_out_533,pxl_out_534,pxl_out_535,pxl_out_536,pxl_out_537,pxl_out_538,pxl_out_539,pxl_out_540,
pxl_out_541,pxl_out_542,pxl_out_543,pxl_out_544,pxl_out_545,pxl_out_546,pxl_out_547,pxl_out_548,pxl_out_549,
pxl_out_550,pxl_out_551,pxl_out_552,pxl_out_553,pxl_out_554,pxl_out_555,pxl_out_556,pxl_out_557,pxl_out_558,
pxl_out_559,pxl_out_560,pxl_out_561,pxl_out_562,pxl_out_563,pxl_out_564,pxl_out_565,pxl_out_566,pxl_out_567,
pxl_out_568,pxl_out_569,pxl_out_570,pxl_out_571,pxl_out_572,pxl_out_573,pxl_out_574,pxl_out_575,pxl_out_576,
pxl_out_577,pxl_out_578,pxl_out_579,pxl_out_580,pxl_out_581,pxl_out_582,pxl_out_583,pxl_out_584,pxl_out_585,
pxl_out_586,pxl_out_587,pxl_out_588,pxl_out_589,pxl_out_590,pxl_out_591,pxl_out_592,pxl_out_593,pxl_out_594,
pxl_out_595,pxl_out_596,pxl_out_597,pxl_out_598,pxl_out_599,pxl_out_600,pxl_out_601,pxl_out_602,pxl_out_603,
pxl_out_604,pxl_out_605,pxl_out_606,pxl_out_607,pxl_out_608,pxl_out_609,pxl_out_610,pxl_out_611,pxl_out_612,
pxl_out_613,pxl_out_614,pxl_out_615,pxl_out_616,pxl_out_617,pxl_out_618,pxl_out_619,pxl_out_620,pxl_out_621,
pxl_out_622,pxl_out_623,pxl_out_624,pxl_out_625,pxl_out_626,pxl_out_627,pxl_out_628,pxl_out_629,pxl_out_630,
pxl_out_631,pxl_out_632,pxl_out_633,pxl_out_634,pxl_out_635,pxl_out_636,pxl_out_637,pxl_out_638,pxl_out_639,
pxl_out_640,pxl_out_641,pxl_out_642,pxl_out_643,pxl_out_644,pxl_out_645,pxl_out_646,pxl_out_647,pxl_out_648,
pxl_out_649,pxl_out_650,pxl_out_651,pxl_out_652,pxl_out_653,pxl_out_654,pxl_out_655,pxl_out_656,pxl_out_657,
pxl_out_658,pxl_out_659,pxl_out_660,pxl_out_661,pxl_out_662,pxl_out_663,pxl_out_664,pxl_out_665,pxl_out_666,
pxl_out_667,pxl_out_668,pxl_out_669,pxl_out_670,pxl_out_671,pxl_out_672,pxl_out_673,pxl_out_674,pxl_out_675,
pxl_out_676,pxl_out_677,pxl_out_678,pxl_out_679,pxl_out_680,pxl_out_681,pxl_out_682,pxl_out_683,pxl_out_684,
pxl_out_685,pxl_out_686,pxl_out_687,pxl_out_688,pxl_out_689,pxl_out_690,pxl_out_691,pxl_out_692,pxl_out_693,
pxl_out_694,pxl_out_695,pxl_out_696,pxl_out_697,pxl_out_698,pxl_out_699,pxl_out_700,pxl_out_701,pxl_out_702,
pxl_out_703,pxl_out_704,pxl_out_705,pxl_out_706,pxl_out_707,pxl_out_708,pxl_out_709,pxl_out_710,pxl_out_711,
pxl_out_712,pxl_out_713,pxl_out_714,pxl_out_715,pxl_out_716,pxl_out_717,pxl_out_718,pxl_out_719,pxl_out_720,
pxl_out_721,pxl_out_722,pxl_out_723,pxl_out_724,pxl_out_725,pxl_out_726,pxl_out_727,pxl_out_728,pxl_out_729,
pxl_out_730,pxl_out_731,pxl_out_732,pxl_out_733,pxl_out_734,pxl_out_735,pxl_out_736,pxl_out_737,pxl_out_738,
pxl_out_739,pxl_out_740,pxl_out_741,pxl_out_742,pxl_out_743,pxl_out_744,pxl_out_745,pxl_out_746,pxl_out_747,
pxl_out_748,pxl_out_749,pxl_out_750,pxl_out_751,pxl_out_752,pxl_out_753,pxl_out_754,pxl_out_755,pxl_out_756,
pxl_out_757,pxl_out_758,pxl_out_759,pxl_out_760,pxl_out_761,pxl_out_762,pxl_out_763,pxl_out_764,pxl_out_765,
pxl_out_766,pxl_out_767,pxl_out_768,pxl_out_769,pxl_out_770,pxl_out_771,pxl_out_772,pxl_out_773,pxl_out_774,
pxl_out_775,pxl_out_776,pxl_out_777,pxl_out_778,pxl_out_779,pxl_out_780,pxl_out_781,pxl_out_782,pxl_out_783,
pxl_out_784,pxl_out_785,pxl_out_786,pxl_out_787,pxl_out_788,pxl_out_789,pxl_out_790,pxl_out_791,pxl_out_792,
pxl_out_793,pxl_out_794,pxl_out_795,pxl_out_796,pxl_out_797,pxl_out_798,pxl_out_799,pxl_out_800,pxl_out_801,
pxl_out_802,pxl_out_803,pxl_out_804,pxl_out_805,pxl_out_806,pxl_out_807,pxl_out_808,pxl_out_809,pxl_out_810,
pxl_out_811,pxl_out_812,pxl_out_813,pxl_out_814,pxl_out_815,pxl_out_816,pxl_out_817,pxl_out_818,pxl_out_819,
pxl_out_820,pxl_out_821,pxl_out_822,pxl_out_823,pxl_out_824,pxl_out_825,pxl_out_826,pxl_out_827,pxl_out_828,
pxl_out_829,pxl_out_830,pxl_out_831,pxl_out_832,pxl_out_833,pxl_out_834,pxl_out_835,pxl_out_836,pxl_out_837,
pxl_out_838,pxl_out_839,pxl_out_840,pxl_out_841,pxl_out_842,pxl_out_843,pxl_out_844,pxl_out_845,pxl_out_846,
pxl_out_847,pxl_out_848,pxl_out_849,pxl_out_850,pxl_out_851,pxl_out_852,pxl_out_853,pxl_out_854,pxl_out_855,
pxl_out_856,pxl_out_857,pxl_out_858,pxl_out_859,pxl_out_860,pxl_out_861,pxl_out_862,pxl_out_863,pxl_out_864,
pxl_out_865,pxl_out_866,pxl_out_867,pxl_out_868,pxl_out_869,pxl_out_870,pxl_out_871,pxl_out_872,pxl_out_873,
pxl_out_874,pxl_out_875,pxl_out_876,pxl_out_877,pxl_out_878,pxl_out_879,pxl_out_880,pxl_out_881,pxl_out_882,
pxl_out_883,pxl_out_884,pxl_out_885,pxl_out_886,pxl_out_887,pxl_out_888,pxl_out_889,pxl_out_890,pxl_out_891,
pxl_out_892,pxl_out_893,pxl_out_894,pxl_out_895,pxl_out_896,pxl_out_897,pxl_out_898,pxl_out_899,pxl_out_900,
pxl_out_901,pxl_out_902,pxl_out_903,pxl_out_904,pxl_out_905,pxl_out_906,pxl_out_907,pxl_out_908,pxl_out_909,
pxl_out_910,pxl_out_911,pxl_out_912,pxl_out_913,pxl_out_914,pxl_out_915,pxl_out_916,pxl_out_917,pxl_out_918,
pxl_out_919,pxl_out_920,pxl_out_921,pxl_out_922,pxl_out_923,pxl_out_924,pxl_out_925,pxl_out_926,pxl_out_927,
pxl_out_928,pxl_out_929,pxl_out_930,pxl_out_931,pxl_out_932,pxl_out_933,pxl_out_934,pxl_out_935,pxl_out_936,
pxl_out_937,pxl_out_938,pxl_out_939,pxl_out_940,pxl_out_941,pxl_out_942,pxl_out_943,pxl_out_944,pxl_out_945,
pxl_out_946,pxl_out_947,pxl_out_948,pxl_out_949,pxl_out_950,pxl_out_951,pxl_out_952,pxl_out_953,pxl_out_954,
pxl_out_955,pxl_out_956,pxl_out_957,pxl_out_958,pxl_out_959,pxl_out_960,pxl_out_961,pxl_out_962,pxl_out_963,
pxl_out_964,pxl_out_965,pxl_out_966,pxl_out_967,pxl_out_968,pxl_out_969,pxl_out_970,pxl_out_971,pxl_out_972,
pxl_out_973,pxl_out_974,pxl_out_975,pxl_out_976,pxl_out_977,pxl_out_978,pxl_out_979,pxl_out_980,pxl_out_981,
pxl_out_982,pxl_out_983,pxl_out_984,pxl_out_985,pxl_out_986,pxl_out_987,pxl_out_988,pxl_out_989,pxl_out_990,
pxl_out_991,pxl_out_992,pxl_out_993,pxl_out_994,pxl_out_995,pxl_out_996,pxl_out_997,pxl_out_998,pxl_out_999,
pxl_out_1000,pxl_out_1001,pxl_out_1002,pxl_out_1003,pxl_out_1004,pxl_out_1005,pxl_out_1006,pxl_out_1007,pxl_out_1008,
pxl_out_1009,pxl_out_1010,pxl_out_1011,pxl_out_1012,pxl_out_1013,pxl_out_1014,pxl_out_1015,pxl_out_1016,pxl_out_1017,
pxl_out_1018,pxl_out_1019,pxl_out_1020,pxl_out_1021,pxl_out_1022,pxl_out_1023,pxl_out_1024;  
  
  wire valid_out_1,valid_out_2,valid_out_3,valid_out_4,valid_out_5,valid_out_6,valid_out_7,valid_out_8,valid_out_9,
valid_out_10,valid_out_11,valid_out_12,valid_out_13,valid_out_14,valid_out_15,valid_out_16,valid_out_17,valid_out_18,
valid_out_19,valid_out_20,valid_out_21,valid_out_22,valid_out_23,valid_out_24,valid_out_25,valid_out_26,valid_out_27,
valid_out_28,valid_out_29,valid_out_30,valid_out_31,valid_out_32,valid_out_33,valid_out_34,valid_out_35,valid_out_36,
valid_out_37,valid_out_38,valid_out_39,valid_out_40,valid_out_41,valid_out_42,valid_out_43,valid_out_44,valid_out_45,
valid_out_46,valid_out_47,valid_out_48,valid_out_49,valid_out_50,valid_out_51,valid_out_52,valid_out_53,valid_out_54,
valid_out_55,valid_out_56,valid_out_57,valid_out_58,valid_out_59,valid_out_60,valid_out_61,valid_out_62,valid_out_63,
valid_out_64,valid_out_65,valid_out_66,valid_out_67,valid_out_68,valid_out_69,valid_out_70,valid_out_71,valid_out_72,
valid_out_73,valid_out_74,valid_out_75,valid_out_76,valid_out_77,valid_out_78,valid_out_79,valid_out_80,valid_out_81,
valid_out_82,valid_out_83,valid_out_84,valid_out_85,valid_out_86,valid_out_87,valid_out_88,valid_out_89,valid_out_90,
valid_out_91,valid_out_92,valid_out_93,valid_out_94,valid_out_95,valid_out_96,valid_out_97,valid_out_98,valid_out_99,
valid_out_100,valid_out_101,valid_out_102,valid_out_103,valid_out_104,valid_out_105,valid_out_106,valid_out_107,valid_out_108,
valid_out_109,valid_out_110,valid_out_111,valid_out_112,valid_out_113,valid_out_114,valid_out_115,valid_out_116,valid_out_117,
valid_out_118,valid_out_119,valid_out_120,valid_out_121,valid_out_122,valid_out_123,valid_out_124,valid_out_125,valid_out_126,
valid_out_127,valid_out_128,valid_out_129,valid_out_130,valid_out_131,valid_out_132,valid_out_133,valid_out_134,valid_out_135,
valid_out_136,valid_out_137,valid_out_138,valid_out_139,valid_out_140,valid_out_141,valid_out_142,valid_out_143,valid_out_144,
valid_out_145,valid_out_146,valid_out_147,valid_out_148,valid_out_149,valid_out_150,valid_out_151,valid_out_152,valid_out_153,
valid_out_154,valid_out_155,valid_out_156,valid_out_157,valid_out_158,valid_out_159,valid_out_160,valid_out_161,valid_out_162,
valid_out_163,valid_out_164,valid_out_165,valid_out_166,valid_out_167,valid_out_168,valid_out_169,valid_out_170,valid_out_171,
valid_out_172,valid_out_173,valid_out_174,valid_out_175,valid_out_176,valid_out_177,valid_out_178,valid_out_179,valid_out_180,
valid_out_181,valid_out_182,valid_out_183,valid_out_184,valid_out_185,valid_out_186,valid_out_187,valid_out_188,valid_out_189,
valid_out_190,valid_out_191,valid_out_192,valid_out_193,valid_out_194,valid_out_195,valid_out_196,valid_out_197,valid_out_198,
valid_out_199,valid_out_200,valid_out_201,valid_out_202,valid_out_203,valid_out_204,valid_out_205,valid_out_206,valid_out_207,
valid_out_208,valid_out_209,valid_out_210,valid_out_211,valid_out_212,valid_out_213,valid_out_214,valid_out_215,valid_out_216,
valid_out_217,valid_out_218,valid_out_219,valid_out_220,valid_out_221,valid_out_222,valid_out_223,valid_out_224,valid_out_225,
valid_out_226,valid_out_227,valid_out_228,valid_out_229,valid_out_230,valid_out_231,valid_out_232,valid_out_233,valid_out_234,
valid_out_235,valid_out_236,valid_out_237,valid_out_238,valid_out_239,valid_out_240,valid_out_241,valid_out_242,valid_out_243,
valid_out_244,valid_out_245,valid_out_246,valid_out_247,valid_out_248,valid_out_249,valid_out_250,valid_out_251,valid_out_252,
valid_out_253,valid_out_254,valid_out_255,valid_out_256,valid_out_257,valid_out_258,valid_out_259,valid_out_260,valid_out_261,
valid_out_262,valid_out_263,valid_out_264,valid_out_265,valid_out_266,valid_out_267,valid_out_268,valid_out_269,valid_out_270,
valid_out_271,valid_out_272,valid_out_273,valid_out_274,valid_out_275,valid_out_276,valid_out_277,valid_out_278,valid_out_279,
valid_out_280,valid_out_281,valid_out_282,valid_out_283,valid_out_284,valid_out_285,valid_out_286,valid_out_287,valid_out_288,
valid_out_289,valid_out_290,valid_out_291,valid_out_292,valid_out_293,valid_out_294,valid_out_295,valid_out_296,valid_out_297,
valid_out_298,valid_out_299,valid_out_300,valid_out_301,valid_out_302,valid_out_303,valid_out_304,valid_out_305,valid_out_306,
valid_out_307,valid_out_308,valid_out_309,valid_out_310,valid_out_311,valid_out_312,valid_out_313,valid_out_314,valid_out_315,
valid_out_316,valid_out_317,valid_out_318,valid_out_319,valid_out_320,valid_out_321,valid_out_322,valid_out_323,valid_out_324,
valid_out_325,valid_out_326,valid_out_327,valid_out_328,valid_out_329,valid_out_330,valid_out_331,valid_out_332,valid_out_333,
valid_out_334,valid_out_335,valid_out_336,valid_out_337,valid_out_338,valid_out_339,valid_out_340,valid_out_341,valid_out_342,
valid_out_343,valid_out_344,valid_out_345,valid_out_346,valid_out_347,valid_out_348,valid_out_349,valid_out_350,valid_out_351,
valid_out_352,valid_out_353,valid_out_354,valid_out_355,valid_out_356,valid_out_357,valid_out_358,valid_out_359,valid_out_360,
valid_out_361,valid_out_362,valid_out_363,valid_out_364,valid_out_365,valid_out_366,valid_out_367,valid_out_368,valid_out_369,
valid_out_370,valid_out_371,valid_out_372,valid_out_373,valid_out_374,valid_out_375,valid_out_376,valid_out_377,valid_out_378,
valid_out_379,valid_out_380,valid_out_381,valid_out_382,valid_out_383,valid_out_384,valid_out_385,valid_out_386,valid_out_387,
valid_out_388,valid_out_389,valid_out_390,valid_out_391,valid_out_392,valid_out_393,valid_out_394,valid_out_395,valid_out_396,
valid_out_397,valid_out_398,valid_out_399,valid_out_400,valid_out_401,valid_out_402,valid_out_403,valid_out_404,valid_out_405,
valid_out_406,valid_out_407,valid_out_408,valid_out_409,valid_out_410,valid_out_411,valid_out_412,valid_out_413,valid_out_414,
valid_out_415,valid_out_416,valid_out_417,valid_out_418,valid_out_419,valid_out_420,valid_out_421,valid_out_422,valid_out_423,
valid_out_424,valid_out_425,valid_out_426,valid_out_427,valid_out_428,valid_out_429,valid_out_430,valid_out_431,valid_out_432,
valid_out_433,valid_out_434,valid_out_435,valid_out_436,valid_out_437,valid_out_438,valid_out_439,valid_out_440,valid_out_441,
valid_out_442,valid_out_443,valid_out_444,valid_out_445,valid_out_446,valid_out_447,valid_out_448,valid_out_449,valid_out_450,
valid_out_451,valid_out_452,valid_out_453,valid_out_454,valid_out_455,valid_out_456,valid_out_457,valid_out_458,valid_out_459,
valid_out_460,valid_out_461,valid_out_462,valid_out_463,valid_out_464,valid_out_465,valid_out_466,valid_out_467,valid_out_468,
valid_out_469,valid_out_470,valid_out_471,valid_out_472,valid_out_473,valid_out_474,valid_out_475,valid_out_476,valid_out_477,
valid_out_478,valid_out_479,valid_out_480,valid_out_481,valid_out_482,valid_out_483,valid_out_484,valid_out_485,valid_out_486,
valid_out_487,valid_out_488,valid_out_489,valid_out_490,valid_out_491,valid_out_492,valid_out_493,valid_out_494,valid_out_495,
valid_out_496,valid_out_497,valid_out_498,valid_out_499,valid_out_500,valid_out_501,valid_out_502,valid_out_503,valid_out_504,
valid_out_505,valid_out_506,valid_out_507,valid_out_508,valid_out_509,valid_out_510,valid_out_511,valid_out_512,valid_out_513,
valid_out_514,valid_out_515,valid_out_516,valid_out_517,valid_out_518,valid_out_519,valid_out_520,valid_out_521,valid_out_522,
valid_out_523,valid_out_524,valid_out_525,valid_out_526,valid_out_527,valid_out_528,valid_out_529,valid_out_530,valid_out_531,
valid_out_532,valid_out_533,valid_out_534,valid_out_535,valid_out_536,valid_out_537,valid_out_538,valid_out_539,valid_out_540,
valid_out_541,valid_out_542,valid_out_543,valid_out_544,valid_out_545,valid_out_546,valid_out_547,valid_out_548,valid_out_549,
valid_out_550,valid_out_551,valid_out_552,valid_out_553,valid_out_554,valid_out_555,valid_out_556,valid_out_557,valid_out_558,
valid_out_559,valid_out_560,valid_out_561,valid_out_562,valid_out_563,valid_out_564,valid_out_565,valid_out_566,valid_out_567,
valid_out_568,valid_out_569,valid_out_570,valid_out_571,valid_out_572,valid_out_573,valid_out_574,valid_out_575,valid_out_576,
valid_out_577,valid_out_578,valid_out_579,valid_out_580,valid_out_581,valid_out_582,valid_out_583,valid_out_584,valid_out_585,
valid_out_586,valid_out_587,valid_out_588,valid_out_589,valid_out_590,valid_out_591,valid_out_592,valid_out_593,valid_out_594,
valid_out_595,valid_out_596,valid_out_597,valid_out_598,valid_out_599,valid_out_600,valid_out_601,valid_out_602,valid_out_603,
valid_out_604,valid_out_605,valid_out_606,valid_out_607,valid_out_608,valid_out_609,valid_out_610,valid_out_611,valid_out_612,
valid_out_613,valid_out_614,valid_out_615,valid_out_616,valid_out_617,valid_out_618,valid_out_619,valid_out_620,valid_out_621,
valid_out_622,valid_out_623,valid_out_624,valid_out_625,valid_out_626,valid_out_627,valid_out_628,valid_out_629,valid_out_630,
valid_out_631,valid_out_632,valid_out_633,valid_out_634,valid_out_635,valid_out_636,valid_out_637,valid_out_638,valid_out_639,
valid_out_640,valid_out_641,valid_out_642,valid_out_643,valid_out_644,valid_out_645,valid_out_646,valid_out_647,valid_out_648,
valid_out_649,valid_out_650,valid_out_651,valid_out_652,valid_out_653,valid_out_654,valid_out_655,valid_out_656,valid_out_657,
valid_out_658,valid_out_659,valid_out_660,valid_out_661,valid_out_662,valid_out_663,valid_out_664,valid_out_665,valid_out_666,
valid_out_667,valid_out_668,valid_out_669,valid_out_670,valid_out_671,valid_out_672,valid_out_673,valid_out_674,valid_out_675,
valid_out_676,valid_out_677,valid_out_678,valid_out_679,valid_out_680,valid_out_681,valid_out_682,valid_out_683,valid_out_684,
valid_out_685,valid_out_686,valid_out_687,valid_out_688,valid_out_689,valid_out_690,valid_out_691,valid_out_692,valid_out_693,
valid_out_694,valid_out_695,valid_out_696,valid_out_697,valid_out_698,valid_out_699,valid_out_700,valid_out_701,valid_out_702,
valid_out_703,valid_out_704,valid_out_705,valid_out_706,valid_out_707,valid_out_708,valid_out_709,valid_out_710,valid_out_711,
valid_out_712,valid_out_713,valid_out_714,valid_out_715,valid_out_716,valid_out_717,valid_out_718,valid_out_719,valid_out_720,
valid_out_721,valid_out_722,valid_out_723,valid_out_724,valid_out_725,valid_out_726,valid_out_727,valid_out_728,valid_out_729,
valid_out_730,valid_out_731,valid_out_732,valid_out_733,valid_out_734,valid_out_735,valid_out_736,valid_out_737,valid_out_738,
valid_out_739,valid_out_740,valid_out_741,valid_out_742,valid_out_743,valid_out_744,valid_out_745,valid_out_746,valid_out_747,
valid_out_748,valid_out_749,valid_out_750,valid_out_751,valid_out_752,valid_out_753,valid_out_754,valid_out_755,valid_out_756,
valid_out_757,valid_out_758,valid_out_759,valid_out_760,valid_out_761,valid_out_762,valid_out_763,valid_out_764,valid_out_765,
valid_out_766,valid_out_767,valid_out_768,valid_out_769,valid_out_770,valid_out_771,valid_out_772,valid_out_773,valid_out_774,
valid_out_775,valid_out_776,valid_out_777,valid_out_778,valid_out_779,valid_out_780,valid_out_781,valid_out_782,valid_out_783,
valid_out_784,valid_out_785,valid_out_786,valid_out_787,valid_out_788,valid_out_789,valid_out_790,valid_out_791,valid_out_792,
valid_out_793,valid_out_794,valid_out_795,valid_out_796,valid_out_797,valid_out_798,valid_out_799,valid_out_800,valid_out_801,
valid_out_802,valid_out_803,valid_out_804,valid_out_805,valid_out_806,valid_out_807,valid_out_808,valid_out_809,valid_out_810,
valid_out_811,valid_out_812,valid_out_813,valid_out_814,valid_out_815,valid_out_816,valid_out_817,valid_out_818,valid_out_819,
valid_out_820,valid_out_821,valid_out_822,valid_out_823,valid_out_824,valid_out_825,valid_out_826,valid_out_827,valid_out_828,
valid_out_829,valid_out_830,valid_out_831,valid_out_832,valid_out_833,valid_out_834,valid_out_835,valid_out_836,valid_out_837,
valid_out_838,valid_out_839,valid_out_840,valid_out_841,valid_out_842,valid_out_843,valid_out_844,valid_out_845,valid_out_846,
valid_out_847,valid_out_848,valid_out_849,valid_out_850,valid_out_851,valid_out_852,valid_out_853,valid_out_854,valid_out_855,
valid_out_856,valid_out_857,valid_out_858,valid_out_859,valid_out_860,valid_out_861,valid_out_862,valid_out_863,valid_out_864,
valid_out_865,valid_out_866,valid_out_867,valid_out_868,valid_out_869,valid_out_870,valid_out_871,valid_out_872,valid_out_873,
valid_out_874,valid_out_875,valid_out_876,valid_out_877,valid_out_878,valid_out_879,valid_out_880,valid_out_881,valid_out_882,
valid_out_883,valid_out_884,valid_out_885,valid_out_886,valid_out_887,valid_out_888,valid_out_889,valid_out_890,valid_out_891,
valid_out_892,valid_out_893,valid_out_894,valid_out_895,valid_out_896,valid_out_897,valid_out_898,valid_out_899,valid_out_900,
valid_out_901,valid_out_902,valid_out_903,valid_out_904,valid_out_905,valid_out_906,valid_out_907,valid_out_908,valid_out_909,
valid_out_910,valid_out_911,valid_out_912,valid_out_913,valid_out_914,valid_out_915,valid_out_916,valid_out_917,valid_out_918,
valid_out_919,valid_out_920,valid_out_921,valid_out_922,valid_out_923,valid_out_924,valid_out_925,valid_out_926,valid_out_927,
valid_out_928,valid_out_929,valid_out_930,valid_out_931,valid_out_932,valid_out_933,valid_out_934,valid_out_935,valid_out_936,
valid_out_937,valid_out_938,valid_out_939,valid_out_940,valid_out_941,valid_out_942,valid_out_943,valid_out_944,valid_out_945,
valid_out_946,valid_out_947,valid_out_948,valid_out_949,valid_out_950,valid_out_951,valid_out_952,valid_out_953,valid_out_954,
valid_out_955,valid_out_956,valid_out_957,valid_out_958,valid_out_959,valid_out_960,valid_out_961,valid_out_962,valid_out_963,
valid_out_964,valid_out_965,valid_out_966,valid_out_967,valid_out_968,valid_out_969,valid_out_970,valid_out_971,valid_out_972,
valid_out_973,valid_out_974,valid_out_975,valid_out_976,valid_out_977,valid_out_978,valid_out_979,valid_out_980,valid_out_981,
valid_out_982,valid_out_983,valid_out_984,valid_out_985,valid_out_986,valid_out_987,valid_out_988,valid_out_989,valid_out_990,
valid_out_991,valid_out_992,valid_out_993,valid_out_994,valid_out_995,valid_out_996,valid_out_997,valid_out_998,valid_out_999,
valid_out_1000,valid_out_1001,valid_out_1002,valid_out_1003,valid_out_1004,valid_out_1005,valid_out_1006,valid_out_1007,valid_out_1008,
valid_out_1009,valid_out_1010,valid_out_1011,valid_out_1012,valid_out_1013,valid_out_1014,valid_out_1015,valid_out_1016,valid_out_1017,
valid_out_1018,valid_out_1019,valid_out_1020,valid_out_1021,valid_out_1022,valid_out_1023,valid_out_1024;
                        
initial begin
 	clk = 0;  
 	i=0;
	reset = 0;

  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In1);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In2);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In3);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In3);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In4);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In5);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In6);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In7);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In8);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In9);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In10);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In11);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In12);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In13);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In14);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In15);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In16);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In17);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In18);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In19);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In20);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In21);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In22);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In23);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In24);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In25);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In26);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In27);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In28);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In29);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In30);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In31);
  $readmemb("E:/Drive/ICDesign_Seminar/Data/ironman_32bit.txt", In32);
  
	end 
	
	always #(C) clk = ~ clk;
	
	always @(posedge clk) begin
	valid_in_1 = 1;
 	valid_in_2 = 1;
 	valid_in_3 = 1;
 	valid_in_4 = 1;
 	valid_in_5 = 1;
 	valid_in_6 = 1;
 	valid_in_7 = 1;
 	valid_in_8 = 1;
 	valid_in_9 = 1;
 	valid_in_10 = 1;
 	valid_in_11 = 1;
 	valid_in_12 = 1;
 	valid_in_13 = 1;
 	valid_in_14 = 1;
 	valid_in_15 = 1;
 	valid_in_16 = 1;
 	valid_in_17 = 1;
 	valid_in_18 = 1;
 	valid_in_19 = 1;
 	valid_in_20 = 1;
 	valid_in_21 = 1;
 	valid_in_22 = 1;
 	valid_in_23 = 1;
 	valid_in_24 = 1;
 	valid_in_25 = 1;
 	valid_in_26 = 1;
 	valid_in_27 = 1;
 	valid_in_28 = 1;
 	valid_in_29 = 1;
 	valid_in_30 = 1;
 	valid_in_31 = 1;
 	valid_in_32 = 1;
 	
  pxl_in_1 = In1[i];
  pxl_in_2 = In2[i];
  pxl_in_3 = In3[i];
  pxl_in_4 = In4[i];
  pxl_in_5 = In5[i];
  pxl_in_6 = In6[i];
  pxl_in_7 = In7[i];
  pxl_in_8 = In8[i];
  pxl_in_9 = In9[i];
  pxl_in_10 = In10[i];
  pxl_in_11 = In11[i];
  pxl_in_12 = In12[i];
  pxl_in_13 = In13[i];
  pxl_in_14 = In14[i];
  pxl_in_15 = In15[i];
  pxl_in_16 = In16[i];
  pxl_in_17 = In17[i];
  pxl_in_18 = In18[i];
  pxl_in_19 = In19[i];
  pxl_in_20 = In20[i];
  pxl_in_21 = In21[i];
  pxl_in_22 = In22[i];
  pxl_in_23 = In23[i];
  pxl_in_24 = In24[i];
  pxl_in_25 = In25[i];
  pxl_in_26 = In26[i];
  pxl_in_27 = In27[i];
  pxl_in_28 = In28[i];
  pxl_in_29 = In29[i];
  pxl_in_30 = In30[i];
  pxl_in_31 = In31[i];
  pxl_in_32 = In32[i];
  #(I) i = i + 1;
  if(i == (T*3)+3) begin
  $finish;
end
end

	Conv2d_2a_3x3_32 #(D,data_width) uut (
		clk, 
		reset, 
            valid_in_1,  valid_in_2,  valid_in_3,  valid_in_4,  valid_in_5,  valid_in_6,
    	       valid_in_7,  valid_in_8,  valid_in_9,  valid_in_10, valid_in_11, valid_in_12,
    	       valid_in_13, valid_in_14, valid_in_15, valid_in_16, valid_in_17, valid_in_18,
    	       valid_in_19, valid_in_20, valid_in_21, valid_in_22, valid_in_23, valid_in_24,
  	         valid_in_25, valid_in_26, valid_in_27, valid_in_28, valid_in_29, valid_in_30,
    	       valid_in_31, valid_in_32,
		
		
		                        pxl_in_1,  pxl_in_2,  pxl_in_3,  pxl_in_4,  pxl_in_5,  pxl_in_6,
    	                       pxl_in_7,  pxl_in_8,  pxl_in_9,  pxl_in_10, pxl_in_11, pxl_in_12,
    	                       pxl_in_13, pxl_in_14, pxl_in_15, pxl_in_16, pxl_in_17, pxl_in_18,
    	                       pxl_in_19, pxl_in_20, pxl_in_21, pxl_in_22, pxl_in_23, pxl_in_24,
    	                       pxl_in_25, pxl_in_26, pxl_in_27, pxl_in_28, pxl_in_29, pxl_in_30,
    	                       pxl_in_31, pxl_in_32,
		
		                    pxl_out_1,pxl_out_2,pxl_out_3,pxl_out_4,pxl_out_5,pxl_out_6,pxl_out_7,pxl_out_8,pxl_out_9,
pxl_out_10,pxl_out_11,pxl_out_12,pxl_out_13,pxl_out_14,pxl_out_15,pxl_out_16,pxl_out_17,pxl_out_18,
pxl_out_19,pxl_out_20,pxl_out_21,pxl_out_22,pxl_out_23,pxl_out_24,pxl_out_25,pxl_out_26,pxl_out_27,
pxl_out_28,pxl_out_29,pxl_out_30,pxl_out_31,pxl_out_32,pxl_out_33,pxl_out_34,pxl_out_35,pxl_out_36,
pxl_out_37,pxl_out_38,pxl_out_39,pxl_out_40,pxl_out_41,pxl_out_42,pxl_out_43,pxl_out_44,pxl_out_45,
pxl_out_46,pxl_out_47,pxl_out_48,pxl_out_49,pxl_out_50,pxl_out_51,pxl_out_52,pxl_out_53,pxl_out_54,
pxl_out_55,pxl_out_56,pxl_out_57,pxl_out_58,pxl_out_59,pxl_out_60,pxl_out_61,pxl_out_62,pxl_out_63,
pxl_out_64,pxl_out_65,pxl_out_66,pxl_out_67,pxl_out_68,pxl_out_69,pxl_out_70,pxl_out_71,pxl_out_72,
pxl_out_73,pxl_out_74,pxl_out_75,pxl_out_76,pxl_out_77,pxl_out_78,pxl_out_79,pxl_out_80,pxl_out_81,
pxl_out_82,pxl_out_83,pxl_out_84,pxl_out_85,pxl_out_86,pxl_out_87,pxl_out_88,pxl_out_89,pxl_out_90,
pxl_out_91,pxl_out_92,pxl_out_93,pxl_out_94,pxl_out_95,pxl_out_96,pxl_out_97,pxl_out_98,pxl_out_99,
pxl_out_100,pxl_out_101,pxl_out_102,pxl_out_103,pxl_out_104,pxl_out_105,pxl_out_106,pxl_out_107,pxl_out_108,
pxl_out_109,pxl_out_110,pxl_out_111,pxl_out_112,pxl_out_113,pxl_out_114,pxl_out_115,pxl_out_116,pxl_out_117,
pxl_out_118,pxl_out_119,pxl_out_120,pxl_out_121,pxl_out_122,pxl_out_123,pxl_out_124,pxl_out_125,pxl_out_126,
pxl_out_127,pxl_out_128,pxl_out_129,pxl_out_130,pxl_out_131,pxl_out_132,pxl_out_133,pxl_out_134,pxl_out_135,
pxl_out_136,pxl_out_137,pxl_out_138,pxl_out_139,pxl_out_140,pxl_out_141,pxl_out_142,pxl_out_143,pxl_out_144,
pxl_out_145,pxl_out_146,pxl_out_147,pxl_out_148,pxl_out_149,pxl_out_150,pxl_out_151,pxl_out_152,pxl_out_153,
pxl_out_154,pxl_out_155,pxl_out_156,pxl_out_157,pxl_out_158,pxl_out_159,pxl_out_160,pxl_out_161,pxl_out_162,
pxl_out_163,pxl_out_164,pxl_out_165,pxl_out_166,pxl_out_167,pxl_out_168,pxl_out_169,pxl_out_170,pxl_out_171,
pxl_out_172,pxl_out_173,pxl_out_174,pxl_out_175,pxl_out_176,pxl_out_177,pxl_out_178,pxl_out_179,pxl_out_180,
pxl_out_181,pxl_out_182,pxl_out_183,pxl_out_184,pxl_out_185,pxl_out_186,pxl_out_187,pxl_out_188,pxl_out_189,
pxl_out_190,pxl_out_191,pxl_out_192,pxl_out_193,pxl_out_194,pxl_out_195,pxl_out_196,pxl_out_197,pxl_out_198,
pxl_out_199,pxl_out_200,pxl_out_201,pxl_out_202,pxl_out_203,pxl_out_204,pxl_out_205,pxl_out_206,pxl_out_207,
pxl_out_208,pxl_out_209,pxl_out_210,pxl_out_211,pxl_out_212,pxl_out_213,pxl_out_214,pxl_out_215,pxl_out_216,
pxl_out_217,pxl_out_218,pxl_out_219,pxl_out_220,pxl_out_221,pxl_out_222,pxl_out_223,pxl_out_224,pxl_out_225,
pxl_out_226,pxl_out_227,pxl_out_228,pxl_out_229,pxl_out_230,pxl_out_231,pxl_out_232,pxl_out_233,pxl_out_234,
pxl_out_235,pxl_out_236,pxl_out_237,pxl_out_238,pxl_out_239,pxl_out_240,pxl_out_241,pxl_out_242,pxl_out_243,
pxl_out_244,pxl_out_245,pxl_out_246,pxl_out_247,pxl_out_248,pxl_out_249,pxl_out_250,pxl_out_251,pxl_out_252,
pxl_out_253,pxl_out_254,pxl_out_255,pxl_out_256,pxl_out_257,pxl_out_258,pxl_out_259,pxl_out_260,pxl_out_261,
pxl_out_262,pxl_out_263,pxl_out_264,pxl_out_265,pxl_out_266,pxl_out_267,pxl_out_268,pxl_out_269,pxl_out_270,
pxl_out_271,pxl_out_272,pxl_out_273,pxl_out_274,pxl_out_275,pxl_out_276,pxl_out_277,pxl_out_278,pxl_out_279,
pxl_out_280,pxl_out_281,pxl_out_282,pxl_out_283,pxl_out_284,pxl_out_285,pxl_out_286,pxl_out_287,pxl_out_288,
pxl_out_289,pxl_out_290,pxl_out_291,pxl_out_292,pxl_out_293,pxl_out_294,pxl_out_295,pxl_out_296,pxl_out_297,
pxl_out_298,pxl_out_299,pxl_out_300,pxl_out_301,pxl_out_302,pxl_out_303,pxl_out_304,pxl_out_305,pxl_out_306,
pxl_out_307,pxl_out_308,pxl_out_309,pxl_out_310,pxl_out_311,pxl_out_312,pxl_out_313,pxl_out_314,pxl_out_315,
pxl_out_316,pxl_out_317,pxl_out_318,pxl_out_319,pxl_out_320,pxl_out_321,pxl_out_322,pxl_out_323,pxl_out_324,
pxl_out_325,pxl_out_326,pxl_out_327,pxl_out_328,pxl_out_329,pxl_out_330,pxl_out_331,pxl_out_332,pxl_out_333,
pxl_out_334,pxl_out_335,pxl_out_336,pxl_out_337,pxl_out_338,pxl_out_339,pxl_out_340,pxl_out_341,pxl_out_342,
pxl_out_343,pxl_out_344,pxl_out_345,pxl_out_346,pxl_out_347,pxl_out_348,pxl_out_349,pxl_out_350,pxl_out_351,
pxl_out_352,pxl_out_353,pxl_out_354,pxl_out_355,pxl_out_356,pxl_out_357,pxl_out_358,pxl_out_359,pxl_out_360,
pxl_out_361,pxl_out_362,pxl_out_363,pxl_out_364,pxl_out_365,pxl_out_366,pxl_out_367,pxl_out_368,pxl_out_369,
pxl_out_370,pxl_out_371,pxl_out_372,pxl_out_373,pxl_out_374,pxl_out_375,pxl_out_376,pxl_out_377,pxl_out_378,
pxl_out_379,pxl_out_380,pxl_out_381,pxl_out_382,pxl_out_383,pxl_out_384,pxl_out_385,pxl_out_386,pxl_out_387,
pxl_out_388,pxl_out_389,pxl_out_390,pxl_out_391,pxl_out_392,pxl_out_393,pxl_out_394,pxl_out_395,pxl_out_396,
pxl_out_397,pxl_out_398,pxl_out_399,pxl_out_400,pxl_out_401,pxl_out_402,pxl_out_403,pxl_out_404,pxl_out_405,
pxl_out_406,pxl_out_407,pxl_out_408,pxl_out_409,pxl_out_410,pxl_out_411,pxl_out_412,pxl_out_413,pxl_out_414,
pxl_out_415,pxl_out_416,pxl_out_417,pxl_out_418,pxl_out_419,pxl_out_420,pxl_out_421,pxl_out_422,pxl_out_423,
pxl_out_424,pxl_out_425,pxl_out_426,pxl_out_427,pxl_out_428,pxl_out_429,pxl_out_430,pxl_out_431,pxl_out_432,
pxl_out_433,pxl_out_434,pxl_out_435,pxl_out_436,pxl_out_437,pxl_out_438,pxl_out_439,pxl_out_440,pxl_out_441,
pxl_out_442,pxl_out_443,pxl_out_444,pxl_out_445,pxl_out_446,pxl_out_447,pxl_out_448,pxl_out_449,pxl_out_450,
pxl_out_451,pxl_out_452,pxl_out_453,pxl_out_454,pxl_out_455,pxl_out_456,pxl_out_457,pxl_out_458,pxl_out_459,
pxl_out_460,pxl_out_461,pxl_out_462,pxl_out_463,pxl_out_464,pxl_out_465,pxl_out_466,pxl_out_467,pxl_out_468,
pxl_out_469,pxl_out_470,pxl_out_471,pxl_out_472,pxl_out_473,pxl_out_474,pxl_out_475,pxl_out_476,pxl_out_477,
pxl_out_478,pxl_out_479,pxl_out_480,pxl_out_481,pxl_out_482,pxl_out_483,pxl_out_484,pxl_out_485,pxl_out_486,
pxl_out_487,pxl_out_488,pxl_out_489,pxl_out_490,pxl_out_491,pxl_out_492,pxl_out_493,pxl_out_494,pxl_out_495,
pxl_out_496,pxl_out_497,pxl_out_498,pxl_out_499,pxl_out_500,pxl_out_501,pxl_out_502,pxl_out_503,pxl_out_504,
pxl_out_505,pxl_out_506,pxl_out_507,pxl_out_508,pxl_out_509,pxl_out_510,pxl_out_511,pxl_out_512,pxl_out_513,
pxl_out_514,pxl_out_515,pxl_out_516,pxl_out_517,pxl_out_518,pxl_out_519,pxl_out_520,pxl_out_521,pxl_out_522,
pxl_out_523,pxl_out_524,pxl_out_525,pxl_out_526,pxl_out_527,pxl_out_528,pxl_out_529,pxl_out_530,pxl_out_531,
pxl_out_532,pxl_out_533,pxl_out_534,pxl_out_535,pxl_out_536,pxl_out_537,pxl_out_538,pxl_out_539,pxl_out_540,
pxl_out_541,pxl_out_542,pxl_out_543,pxl_out_544,pxl_out_545,pxl_out_546,pxl_out_547,pxl_out_548,pxl_out_549,
pxl_out_550,pxl_out_551,pxl_out_552,pxl_out_553,pxl_out_554,pxl_out_555,pxl_out_556,pxl_out_557,pxl_out_558,
pxl_out_559,pxl_out_560,pxl_out_561,pxl_out_562,pxl_out_563,pxl_out_564,pxl_out_565,pxl_out_566,pxl_out_567,
pxl_out_568,pxl_out_569,pxl_out_570,pxl_out_571,pxl_out_572,pxl_out_573,pxl_out_574,pxl_out_575,pxl_out_576,
pxl_out_577,pxl_out_578,pxl_out_579,pxl_out_580,pxl_out_581,pxl_out_582,pxl_out_583,pxl_out_584,pxl_out_585,
pxl_out_586,pxl_out_587,pxl_out_588,pxl_out_589,pxl_out_590,pxl_out_591,pxl_out_592,pxl_out_593,pxl_out_594,
pxl_out_595,pxl_out_596,pxl_out_597,pxl_out_598,pxl_out_599,pxl_out_600,pxl_out_601,pxl_out_602,pxl_out_603,
pxl_out_604,pxl_out_605,pxl_out_606,pxl_out_607,pxl_out_608,pxl_out_609,pxl_out_610,pxl_out_611,pxl_out_612,
pxl_out_613,pxl_out_614,pxl_out_615,pxl_out_616,pxl_out_617,pxl_out_618,pxl_out_619,pxl_out_620,pxl_out_621,
pxl_out_622,pxl_out_623,pxl_out_624,pxl_out_625,pxl_out_626,pxl_out_627,pxl_out_628,pxl_out_629,pxl_out_630,
pxl_out_631,pxl_out_632,pxl_out_633,pxl_out_634,pxl_out_635,pxl_out_636,pxl_out_637,pxl_out_638,pxl_out_639,
pxl_out_640,pxl_out_641,pxl_out_642,pxl_out_643,pxl_out_644,pxl_out_645,pxl_out_646,pxl_out_647,pxl_out_648,
pxl_out_649,pxl_out_650,pxl_out_651,pxl_out_652,pxl_out_653,pxl_out_654,pxl_out_655,pxl_out_656,pxl_out_657,
pxl_out_658,pxl_out_659,pxl_out_660,pxl_out_661,pxl_out_662,pxl_out_663,pxl_out_664,pxl_out_665,pxl_out_666,
pxl_out_667,pxl_out_668,pxl_out_669,pxl_out_670,pxl_out_671,pxl_out_672,pxl_out_673,pxl_out_674,pxl_out_675,
pxl_out_676,pxl_out_677,pxl_out_678,pxl_out_679,pxl_out_680,pxl_out_681,pxl_out_682,pxl_out_683,pxl_out_684,
pxl_out_685,pxl_out_686,pxl_out_687,pxl_out_688,pxl_out_689,pxl_out_690,pxl_out_691,pxl_out_692,pxl_out_693,
pxl_out_694,pxl_out_695,pxl_out_696,pxl_out_697,pxl_out_698,pxl_out_699,pxl_out_700,pxl_out_701,pxl_out_702,
pxl_out_703,pxl_out_704,pxl_out_705,pxl_out_706,pxl_out_707,pxl_out_708,pxl_out_709,pxl_out_710,pxl_out_711,
pxl_out_712,pxl_out_713,pxl_out_714,pxl_out_715,pxl_out_716,pxl_out_717,pxl_out_718,pxl_out_719,pxl_out_720,
pxl_out_721,pxl_out_722,pxl_out_723,pxl_out_724,pxl_out_725,pxl_out_726,pxl_out_727,pxl_out_728,pxl_out_729,
pxl_out_730,pxl_out_731,pxl_out_732,pxl_out_733,pxl_out_734,pxl_out_735,pxl_out_736,pxl_out_737,pxl_out_738,
pxl_out_739,pxl_out_740,pxl_out_741,pxl_out_742,pxl_out_743,pxl_out_744,pxl_out_745,pxl_out_746,pxl_out_747,
pxl_out_748,pxl_out_749,pxl_out_750,pxl_out_751,pxl_out_752,pxl_out_753,pxl_out_754,pxl_out_755,pxl_out_756,
pxl_out_757,pxl_out_758,pxl_out_759,pxl_out_760,pxl_out_761,pxl_out_762,pxl_out_763,pxl_out_764,pxl_out_765,
pxl_out_766,pxl_out_767,pxl_out_768,pxl_out_769,pxl_out_770,pxl_out_771,pxl_out_772,pxl_out_773,pxl_out_774,
pxl_out_775,pxl_out_776,pxl_out_777,pxl_out_778,pxl_out_779,pxl_out_780,pxl_out_781,pxl_out_782,pxl_out_783,
pxl_out_784,pxl_out_785,pxl_out_786,pxl_out_787,pxl_out_788,pxl_out_789,pxl_out_790,pxl_out_791,pxl_out_792,
pxl_out_793,pxl_out_794,pxl_out_795,pxl_out_796,pxl_out_797,pxl_out_798,pxl_out_799,pxl_out_800,pxl_out_801,
pxl_out_802,pxl_out_803,pxl_out_804,pxl_out_805,pxl_out_806,pxl_out_807,pxl_out_808,pxl_out_809,pxl_out_810,
pxl_out_811,pxl_out_812,pxl_out_813,pxl_out_814,pxl_out_815,pxl_out_816,pxl_out_817,pxl_out_818,pxl_out_819,
pxl_out_820,pxl_out_821,pxl_out_822,pxl_out_823,pxl_out_824,pxl_out_825,pxl_out_826,pxl_out_827,pxl_out_828,
pxl_out_829,pxl_out_830,pxl_out_831,pxl_out_832,pxl_out_833,pxl_out_834,pxl_out_835,pxl_out_836,pxl_out_837,
pxl_out_838,pxl_out_839,pxl_out_840,pxl_out_841,pxl_out_842,pxl_out_843,pxl_out_844,pxl_out_845,pxl_out_846,
pxl_out_847,pxl_out_848,pxl_out_849,pxl_out_850,pxl_out_851,pxl_out_852,pxl_out_853,pxl_out_854,pxl_out_855,
pxl_out_856,pxl_out_857,pxl_out_858,pxl_out_859,pxl_out_860,pxl_out_861,pxl_out_862,pxl_out_863,pxl_out_864,
pxl_out_865,pxl_out_866,pxl_out_867,pxl_out_868,pxl_out_869,pxl_out_870,pxl_out_871,pxl_out_872,pxl_out_873,
pxl_out_874,pxl_out_875,pxl_out_876,pxl_out_877,pxl_out_878,pxl_out_879,pxl_out_880,pxl_out_881,pxl_out_882,
pxl_out_883,pxl_out_884,pxl_out_885,pxl_out_886,pxl_out_887,pxl_out_888,pxl_out_889,pxl_out_890,pxl_out_891,
pxl_out_892,pxl_out_893,pxl_out_894,pxl_out_895,pxl_out_896,pxl_out_897,pxl_out_898,pxl_out_899,pxl_out_900,
pxl_out_901,pxl_out_902,pxl_out_903,pxl_out_904,pxl_out_905,pxl_out_906,pxl_out_907,pxl_out_908,pxl_out_909,
pxl_out_910,pxl_out_911,pxl_out_912,pxl_out_913,pxl_out_914,pxl_out_915,pxl_out_916,pxl_out_917,pxl_out_918,
pxl_out_919,pxl_out_920,pxl_out_921,pxl_out_922,pxl_out_923,pxl_out_924,pxl_out_925,pxl_out_926,pxl_out_927,
pxl_out_928,pxl_out_929,pxl_out_930,pxl_out_931,pxl_out_932,pxl_out_933,pxl_out_934,pxl_out_935,pxl_out_936,
pxl_out_937,pxl_out_938,pxl_out_939,pxl_out_940,pxl_out_941,pxl_out_942,pxl_out_943,pxl_out_944,pxl_out_945,
pxl_out_946,pxl_out_947,pxl_out_948,pxl_out_949,pxl_out_950,pxl_out_951,pxl_out_952,pxl_out_953,pxl_out_954,
pxl_out_955,pxl_out_956,pxl_out_957,pxl_out_958,pxl_out_959,pxl_out_960,pxl_out_961,pxl_out_962,pxl_out_963,
pxl_out_964,pxl_out_965,pxl_out_966,pxl_out_967,pxl_out_968,pxl_out_969,pxl_out_970,pxl_out_971,pxl_out_972,
pxl_out_973,pxl_out_974,pxl_out_975,pxl_out_976,pxl_out_977,pxl_out_978,pxl_out_979,pxl_out_980,pxl_out_981,
pxl_out_982,pxl_out_983,pxl_out_984,pxl_out_985,pxl_out_986,pxl_out_987,pxl_out_988,pxl_out_989,pxl_out_990,
pxl_out_991,pxl_out_992,pxl_out_993,pxl_out_994,pxl_out_995,pxl_out_996,pxl_out_997,pxl_out_998,pxl_out_999,
pxl_out_1000,pxl_out_1001,pxl_out_1002,pxl_out_1003,pxl_out_1004,pxl_out_1005,pxl_out_1006,pxl_out_1007,pxl_out_1008,
pxl_out_1009,pxl_out_1010,pxl_out_1011,pxl_out_1012,pxl_out_1013,pxl_out_1014,pxl_out_1015,pxl_out_1016,pxl_out_1017,
pxl_out_1018,pxl_out_1019,pxl_out_1020,pxl_out_1021,pxl_out_1022,pxl_out_1023,pxl_out_1024,  
  
   valid_out_1,valid_out_2,valid_out_3,valid_out_4,valid_out_5,valid_out_6,valid_out_7,valid_out_8,valid_out_9,
valid_out_10,valid_out_11,valid_out_12,valid_out_13,valid_out_14,valid_out_15,valid_out_16,valid_out_17,valid_out_18,
valid_out_19,valid_out_20,valid_out_21,valid_out_22,valid_out_23,valid_out_24,valid_out_25,valid_out_26,valid_out_27,
valid_out_28,valid_out_29,valid_out_30,valid_out_31,valid_out_32,valid_out_33,valid_out_34,valid_out_35,valid_out_36,
valid_out_37,valid_out_38,valid_out_39,valid_out_40,valid_out_41,valid_out_42,valid_out_43,valid_out_44,valid_out_45,
valid_out_46,valid_out_47,valid_out_48,valid_out_49,valid_out_50,valid_out_51,valid_out_52,valid_out_53,valid_out_54,
valid_out_55,valid_out_56,valid_out_57,valid_out_58,valid_out_59,valid_out_60,valid_out_61,valid_out_62,valid_out_63,
valid_out_64,valid_out_65,valid_out_66,valid_out_67,valid_out_68,valid_out_69,valid_out_70,valid_out_71,valid_out_72,
valid_out_73,valid_out_74,valid_out_75,valid_out_76,valid_out_77,valid_out_78,valid_out_79,valid_out_80,valid_out_81,
valid_out_82,valid_out_83,valid_out_84,valid_out_85,valid_out_86,valid_out_87,valid_out_88,valid_out_89,valid_out_90,
valid_out_91,valid_out_92,valid_out_93,valid_out_94,valid_out_95,valid_out_96,valid_out_97,valid_out_98,valid_out_99,
valid_out_100,valid_out_101,valid_out_102,valid_out_103,valid_out_104,valid_out_105,valid_out_106,valid_out_107,valid_out_108,
valid_out_109,valid_out_110,valid_out_111,valid_out_112,valid_out_113,valid_out_114,valid_out_115,valid_out_116,valid_out_117,
valid_out_118,valid_out_119,valid_out_120,valid_out_121,valid_out_122,valid_out_123,valid_out_124,valid_out_125,valid_out_126,
valid_out_127,valid_out_128,valid_out_129,valid_out_130,valid_out_131,valid_out_132,valid_out_133,valid_out_134,valid_out_135,
valid_out_136,valid_out_137,valid_out_138,valid_out_139,valid_out_140,valid_out_141,valid_out_142,valid_out_143,valid_out_144,
valid_out_145,valid_out_146,valid_out_147,valid_out_148,valid_out_149,valid_out_150,valid_out_151,valid_out_152,valid_out_153,
valid_out_154,valid_out_155,valid_out_156,valid_out_157,valid_out_158,valid_out_159,valid_out_160,valid_out_161,valid_out_162,
valid_out_163,valid_out_164,valid_out_165,valid_out_166,valid_out_167,valid_out_168,valid_out_169,valid_out_170,valid_out_171,
valid_out_172,valid_out_173,valid_out_174,valid_out_175,valid_out_176,valid_out_177,valid_out_178,valid_out_179,valid_out_180,
valid_out_181,valid_out_182,valid_out_183,valid_out_184,valid_out_185,valid_out_186,valid_out_187,valid_out_188,valid_out_189,
valid_out_190,valid_out_191,valid_out_192,valid_out_193,valid_out_194,valid_out_195,valid_out_196,valid_out_197,valid_out_198,
valid_out_199,valid_out_200,valid_out_201,valid_out_202,valid_out_203,valid_out_204,valid_out_205,valid_out_206,valid_out_207,
valid_out_208,valid_out_209,valid_out_210,valid_out_211,valid_out_212,valid_out_213,valid_out_214,valid_out_215,valid_out_216,
valid_out_217,valid_out_218,valid_out_219,valid_out_220,valid_out_221,valid_out_222,valid_out_223,valid_out_224,valid_out_225,
valid_out_226,valid_out_227,valid_out_228,valid_out_229,valid_out_230,valid_out_231,valid_out_232,valid_out_233,valid_out_234,
valid_out_235,valid_out_236,valid_out_237,valid_out_238,valid_out_239,valid_out_240,valid_out_241,valid_out_242,valid_out_243,
valid_out_244,valid_out_245,valid_out_246,valid_out_247,valid_out_248,valid_out_249,valid_out_250,valid_out_251,valid_out_252,
valid_out_253,valid_out_254,valid_out_255,valid_out_256,valid_out_257,valid_out_258,valid_out_259,valid_out_260,valid_out_261,
valid_out_262,valid_out_263,valid_out_264,valid_out_265,valid_out_266,valid_out_267,valid_out_268,valid_out_269,valid_out_270,
valid_out_271,valid_out_272,valid_out_273,valid_out_274,valid_out_275,valid_out_276,valid_out_277,valid_out_278,valid_out_279,
valid_out_280,valid_out_281,valid_out_282,valid_out_283,valid_out_284,valid_out_285,valid_out_286,valid_out_287,valid_out_288,
valid_out_289,valid_out_290,valid_out_291,valid_out_292,valid_out_293,valid_out_294,valid_out_295,valid_out_296,valid_out_297,
valid_out_298,valid_out_299,valid_out_300,valid_out_301,valid_out_302,valid_out_303,valid_out_304,valid_out_305,valid_out_306,
valid_out_307,valid_out_308,valid_out_309,valid_out_310,valid_out_311,valid_out_312,valid_out_313,valid_out_314,valid_out_315,
valid_out_316,valid_out_317,valid_out_318,valid_out_319,valid_out_320,valid_out_321,valid_out_322,valid_out_323,valid_out_324,
valid_out_325,valid_out_326,valid_out_327,valid_out_328,valid_out_329,valid_out_330,valid_out_331,valid_out_332,valid_out_333,
valid_out_334,valid_out_335,valid_out_336,valid_out_337,valid_out_338,valid_out_339,valid_out_340,valid_out_341,valid_out_342,
valid_out_343,valid_out_344,valid_out_345,valid_out_346,valid_out_347,valid_out_348,valid_out_349,valid_out_350,valid_out_351,
valid_out_352,valid_out_353,valid_out_354,valid_out_355,valid_out_356,valid_out_357,valid_out_358,valid_out_359,valid_out_360,
valid_out_361,valid_out_362,valid_out_363,valid_out_364,valid_out_365,valid_out_366,valid_out_367,valid_out_368,valid_out_369,
valid_out_370,valid_out_371,valid_out_372,valid_out_373,valid_out_374,valid_out_375,valid_out_376,valid_out_377,valid_out_378,
valid_out_379,valid_out_380,valid_out_381,valid_out_382,valid_out_383,valid_out_384,valid_out_385,valid_out_386,valid_out_387,
valid_out_388,valid_out_389,valid_out_390,valid_out_391,valid_out_392,valid_out_393,valid_out_394,valid_out_395,valid_out_396,
valid_out_397,valid_out_398,valid_out_399,valid_out_400,valid_out_401,valid_out_402,valid_out_403,valid_out_404,valid_out_405,
valid_out_406,valid_out_407,valid_out_408,valid_out_409,valid_out_410,valid_out_411,valid_out_412,valid_out_413,valid_out_414,
valid_out_415,valid_out_416,valid_out_417,valid_out_418,valid_out_419,valid_out_420,valid_out_421,valid_out_422,valid_out_423,
valid_out_424,valid_out_425,valid_out_426,valid_out_427,valid_out_428,valid_out_429,valid_out_430,valid_out_431,valid_out_432,
valid_out_433,valid_out_434,valid_out_435,valid_out_436,valid_out_437,valid_out_438,valid_out_439,valid_out_440,valid_out_441,
valid_out_442,valid_out_443,valid_out_444,valid_out_445,valid_out_446,valid_out_447,valid_out_448,valid_out_449,valid_out_450,
valid_out_451,valid_out_452,valid_out_453,valid_out_454,valid_out_455,valid_out_456,valid_out_457,valid_out_458,valid_out_459,
valid_out_460,valid_out_461,valid_out_462,valid_out_463,valid_out_464,valid_out_465,valid_out_466,valid_out_467,valid_out_468,
valid_out_469,valid_out_470,valid_out_471,valid_out_472,valid_out_473,valid_out_474,valid_out_475,valid_out_476,valid_out_477,
valid_out_478,valid_out_479,valid_out_480,valid_out_481,valid_out_482,valid_out_483,valid_out_484,valid_out_485,valid_out_486,
valid_out_487,valid_out_488,valid_out_489,valid_out_490,valid_out_491,valid_out_492,valid_out_493,valid_out_494,valid_out_495,
valid_out_496,valid_out_497,valid_out_498,valid_out_499,valid_out_500,valid_out_501,valid_out_502,valid_out_503,valid_out_504,
valid_out_505,valid_out_506,valid_out_507,valid_out_508,valid_out_509,valid_out_510,valid_out_511,valid_out_512,valid_out_513,
valid_out_514,valid_out_515,valid_out_516,valid_out_517,valid_out_518,valid_out_519,valid_out_520,valid_out_521,valid_out_522,
valid_out_523,valid_out_524,valid_out_525,valid_out_526,valid_out_527,valid_out_528,valid_out_529,valid_out_530,valid_out_531,
valid_out_532,valid_out_533,valid_out_534,valid_out_535,valid_out_536,valid_out_537,valid_out_538,valid_out_539,valid_out_540,
valid_out_541,valid_out_542,valid_out_543,valid_out_544,valid_out_545,valid_out_546,valid_out_547,valid_out_548,valid_out_549,
valid_out_550,valid_out_551,valid_out_552,valid_out_553,valid_out_554,valid_out_555,valid_out_556,valid_out_557,valid_out_558,
valid_out_559,valid_out_560,valid_out_561,valid_out_562,valid_out_563,valid_out_564,valid_out_565,valid_out_566,valid_out_567,
valid_out_568,valid_out_569,valid_out_570,valid_out_571,valid_out_572,valid_out_573,valid_out_574,valid_out_575,valid_out_576,
valid_out_577,valid_out_578,valid_out_579,valid_out_580,valid_out_581,valid_out_582,valid_out_583,valid_out_584,valid_out_585,
valid_out_586,valid_out_587,valid_out_588,valid_out_589,valid_out_590,valid_out_591,valid_out_592,valid_out_593,valid_out_594,
valid_out_595,valid_out_596,valid_out_597,valid_out_598,valid_out_599,valid_out_600,valid_out_601,valid_out_602,valid_out_603,
valid_out_604,valid_out_605,valid_out_606,valid_out_607,valid_out_608,valid_out_609,valid_out_610,valid_out_611,valid_out_612,
valid_out_613,valid_out_614,valid_out_615,valid_out_616,valid_out_617,valid_out_618,valid_out_619,valid_out_620,valid_out_621,
valid_out_622,valid_out_623,valid_out_624,valid_out_625,valid_out_626,valid_out_627,valid_out_628,valid_out_629,valid_out_630,
valid_out_631,valid_out_632,valid_out_633,valid_out_634,valid_out_635,valid_out_636,valid_out_637,valid_out_638,valid_out_639,
valid_out_640,valid_out_641,valid_out_642,valid_out_643,valid_out_644,valid_out_645,valid_out_646,valid_out_647,valid_out_648,
valid_out_649,valid_out_650,valid_out_651,valid_out_652,valid_out_653,valid_out_654,valid_out_655,valid_out_656,valid_out_657,
valid_out_658,valid_out_659,valid_out_660,valid_out_661,valid_out_662,valid_out_663,valid_out_664,valid_out_665,valid_out_666,
valid_out_667,valid_out_668,valid_out_669,valid_out_670,valid_out_671,valid_out_672,valid_out_673,valid_out_674,valid_out_675,
valid_out_676,valid_out_677,valid_out_678,valid_out_679,valid_out_680,valid_out_681,valid_out_682,valid_out_683,valid_out_684,
valid_out_685,valid_out_686,valid_out_687,valid_out_688,valid_out_689,valid_out_690,valid_out_691,valid_out_692,valid_out_693,
valid_out_694,valid_out_695,valid_out_696,valid_out_697,valid_out_698,valid_out_699,valid_out_700,valid_out_701,valid_out_702,
valid_out_703,valid_out_704,valid_out_705,valid_out_706,valid_out_707,valid_out_708,valid_out_709,valid_out_710,valid_out_711,
valid_out_712,valid_out_713,valid_out_714,valid_out_715,valid_out_716,valid_out_717,valid_out_718,valid_out_719,valid_out_720,
valid_out_721,valid_out_722,valid_out_723,valid_out_724,valid_out_725,valid_out_726,valid_out_727,valid_out_728,valid_out_729,
valid_out_730,valid_out_731,valid_out_732,valid_out_733,valid_out_734,valid_out_735,valid_out_736,valid_out_737,valid_out_738,
valid_out_739,valid_out_740,valid_out_741,valid_out_742,valid_out_743,valid_out_744,valid_out_745,valid_out_746,valid_out_747,
valid_out_748,valid_out_749,valid_out_750,valid_out_751,valid_out_752,valid_out_753,valid_out_754,valid_out_755,valid_out_756,
valid_out_757,valid_out_758,valid_out_759,valid_out_760,valid_out_761,valid_out_762,valid_out_763,valid_out_764,valid_out_765,
valid_out_766,valid_out_767,valid_out_768,valid_out_769,valid_out_770,valid_out_771,valid_out_772,valid_out_773,valid_out_774,
valid_out_775,valid_out_776,valid_out_777,valid_out_778,valid_out_779,valid_out_780,valid_out_781,valid_out_782,valid_out_783,
valid_out_784,valid_out_785,valid_out_786,valid_out_787,valid_out_788,valid_out_789,valid_out_790,valid_out_791,valid_out_792,
valid_out_793,valid_out_794,valid_out_795,valid_out_796,valid_out_797,valid_out_798,valid_out_799,valid_out_800,valid_out_801,
valid_out_802,valid_out_803,valid_out_804,valid_out_805,valid_out_806,valid_out_807,valid_out_808,valid_out_809,valid_out_810,
valid_out_811,valid_out_812,valid_out_813,valid_out_814,valid_out_815,valid_out_816,valid_out_817,valid_out_818,valid_out_819,
valid_out_820,valid_out_821,valid_out_822,valid_out_823,valid_out_824,valid_out_825,valid_out_826,valid_out_827,valid_out_828,
valid_out_829,valid_out_830,valid_out_831,valid_out_832,valid_out_833,valid_out_834,valid_out_835,valid_out_836,valid_out_837,
valid_out_838,valid_out_839,valid_out_840,valid_out_841,valid_out_842,valid_out_843,valid_out_844,valid_out_845,valid_out_846,
valid_out_847,valid_out_848,valid_out_849,valid_out_850,valid_out_851,valid_out_852,valid_out_853,valid_out_854,valid_out_855,
valid_out_856,valid_out_857,valid_out_858,valid_out_859,valid_out_860,valid_out_861,valid_out_862,valid_out_863,valid_out_864,
valid_out_865,valid_out_866,valid_out_867,valid_out_868,valid_out_869,valid_out_870,valid_out_871,valid_out_872,valid_out_873,
valid_out_874,valid_out_875,valid_out_876,valid_out_877,valid_out_878,valid_out_879,valid_out_880,valid_out_881,valid_out_882,
valid_out_883,valid_out_884,valid_out_885,valid_out_886,valid_out_887,valid_out_888,valid_out_889,valid_out_890,valid_out_891,
valid_out_892,valid_out_893,valid_out_894,valid_out_895,valid_out_896,valid_out_897,valid_out_898,valid_out_899,valid_out_900,
valid_out_901,valid_out_902,valid_out_903,valid_out_904,valid_out_905,valid_out_906,valid_out_907,valid_out_908,valid_out_909,
valid_out_910,valid_out_911,valid_out_912,valid_out_913,valid_out_914,valid_out_915,valid_out_916,valid_out_917,valid_out_918,
valid_out_919,valid_out_920,valid_out_921,valid_out_922,valid_out_923,valid_out_924,valid_out_925,valid_out_926,valid_out_927,
valid_out_928,valid_out_929,valid_out_930,valid_out_931,valid_out_932,valid_out_933,valid_out_934,valid_out_935,valid_out_936,
valid_out_937,valid_out_938,valid_out_939,valid_out_940,valid_out_941,valid_out_942,valid_out_943,valid_out_944,valid_out_945,
valid_out_946,valid_out_947,valid_out_948,valid_out_949,valid_out_950,valid_out_951,valid_out_952,valid_out_953,valid_out_954,
valid_out_955,valid_out_956,valid_out_957,valid_out_958,valid_out_959,valid_out_960,valid_out_961,valid_out_962,valid_out_963,
valid_out_964,valid_out_965,valid_out_966,valid_out_967,valid_out_968,valid_out_969,valid_out_970,valid_out_971,valid_out_972,
valid_out_973,valid_out_974,valid_out_975,valid_out_976,valid_out_977,valid_out_978,valid_out_979,valid_out_980,valid_out_981,
valid_out_982,valid_out_983,valid_out_984,valid_out_985,valid_out_986,valid_out_987,valid_out_988,valid_out_989,valid_out_990,
valid_out_991,valid_out_992,valid_out_993,valid_out_994,valid_out_995,valid_out_996,valid_out_997,valid_out_998,valid_out_999,
valid_out_1000,valid_out_1001,valid_out_1002,valid_out_1003,valid_out_1004,valid_out_1005,valid_out_1006,valid_out_1007,valid_out_1008,
valid_out_1009,valid_out_1010,valid_out_1011,valid_out_1012,valid_out_1013,valid_out_1014,valid_out_1015,valid_out_1016,valid_out_1017,
valid_out_1018,valid_out_1019,valid_out_1020,valid_out_1021,valid_out_1022,valid_out_1023,valid_out_1024  

	);

endmodule                      

