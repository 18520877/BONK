// add 3 input to 1 input
// 147x147x1024 -> 147x147x32

 module add_1024to32
#(
  parameter D = 220,
  parameter DATA_WIDTH = 32)
(
    	input clk,
     	input reset,
     	input valid_in_1,valid_in_2,valid_in_3,valid_in_4,valid_in_5,valid_in_6,valid_in_7,valid_in_8,valid_in_9,
valid_in_10,valid_in_11,valid_in_12,valid_in_13,valid_in_14,valid_in_15,valid_in_16,valid_in_17,valid_in_18,
valid_in_19,valid_in_20,valid_in_21,valid_in_22,valid_in_23,valid_in_24,valid_in_25,valid_in_26,valid_in_27,
valid_in_28,valid_in_29,valid_in_30,valid_in_31,valid_in_32,valid_in_33,valid_in_34,valid_in_35,valid_in_36,
valid_in_37,valid_in_38,valid_in_39,valid_in_40,valid_in_41,valid_in_42,valid_in_43,valid_in_44,valid_in_45,
valid_in_46,valid_in_47,valid_in_48,valid_in_49,valid_in_50,valid_in_51,valid_in_52,valid_in_53,valid_in_54,
valid_in_55,valid_in_56,valid_in_57,valid_in_58,valid_in_59,valid_in_60,valid_in_61,valid_in_62,valid_in_63,
valid_in_64,valid_in_65,valid_in_66,valid_in_67,valid_in_68,valid_in_69,valid_in_70,valid_in_71,valid_in_72,
valid_in_73,valid_in_74,valid_in_75,valid_in_76,valid_in_77,valid_in_78,valid_in_79,valid_in_80,valid_in_81,
valid_in_82,valid_in_83,valid_in_84,valid_in_85,valid_in_86,valid_in_87,valid_in_88,valid_in_89,valid_in_90,
valid_in_91,valid_in_92,valid_in_93,valid_in_94,valid_in_95,valid_in_96,valid_in_97,valid_in_98,valid_in_99,
valid_in_100,valid_in_101,valid_in_102,valid_in_103,valid_in_104,valid_in_105,valid_in_106,valid_in_107,valid_in_108,
valid_in_109,valid_in_110,valid_in_111,valid_in_112,valid_in_113,valid_in_114,valid_in_115,valid_in_116,valid_in_117,
valid_in_118,valid_in_119,valid_in_120,valid_in_121,valid_in_122,valid_in_123,valid_in_124,valid_in_125,valid_in_126,
valid_in_127,valid_in_128,valid_in_129,valid_in_130,valid_in_131,valid_in_132,valid_in_133,valid_in_134,valid_in_135,
valid_in_136,valid_in_137,valid_in_138,valid_in_139,valid_in_140,valid_in_141,valid_in_142,valid_in_143,valid_in_144,
valid_in_145,valid_in_146,valid_in_147,valid_in_148,valid_in_149,valid_in_150,valid_in_151,valid_in_152,valid_in_153,
valid_in_154,valid_in_155,valid_in_156,valid_in_157,valid_in_158,valid_in_159,valid_in_160,valid_in_161,valid_in_162,
valid_in_163,valid_in_164,valid_in_165,valid_in_166,valid_in_167,valid_in_168,valid_in_169,valid_in_170,valid_in_171,
valid_in_172,valid_in_173,valid_in_174,valid_in_175,valid_in_176,valid_in_177,valid_in_178,valid_in_179,valid_in_180,
valid_in_181,valid_in_182,valid_in_183,valid_in_184,valid_in_185,valid_in_186,valid_in_187,valid_in_188,valid_in_189,
valid_in_190,valid_in_191,valid_in_192,valid_in_193,valid_in_194,valid_in_195,valid_in_196,valid_in_197,valid_in_198,
valid_in_199,valid_in_200,valid_in_201,valid_in_202,valid_in_203,valid_in_204,valid_in_205,valid_in_206,valid_in_207,
valid_in_208,valid_in_209,valid_in_210,valid_in_211,valid_in_212,valid_in_213,valid_in_214,valid_in_215,valid_in_216,
valid_in_217,valid_in_218,valid_in_219,valid_in_220,valid_in_221,valid_in_222,valid_in_223,valid_in_224,valid_in_225,
valid_in_226,valid_in_227,valid_in_228,valid_in_229,valid_in_230,valid_in_231,valid_in_232,valid_in_233,valid_in_234,
valid_in_235,valid_in_236,valid_in_237,valid_in_238,valid_in_239,valid_in_240,valid_in_241,valid_in_242,valid_in_243,
valid_in_244,valid_in_245,valid_in_246,valid_in_247,valid_in_248,valid_in_249,valid_in_250,valid_in_251,valid_in_252,
valid_in_253,valid_in_254,valid_in_255,valid_in_256,valid_in_257,valid_in_258,valid_in_259,valid_in_260,valid_in_261,
valid_in_262,valid_in_263,valid_in_264,valid_in_265,valid_in_266,valid_in_267,valid_in_268,valid_in_269,valid_in_270,
valid_in_271,valid_in_272,valid_in_273,valid_in_274,valid_in_275,valid_in_276,valid_in_277,valid_in_278,valid_in_279,
valid_in_280,valid_in_281,valid_in_282,valid_in_283,valid_in_284,valid_in_285,valid_in_286,valid_in_287,valid_in_288,
valid_in_289,valid_in_290,valid_in_291,valid_in_292,valid_in_293,valid_in_294,valid_in_295,valid_in_296,valid_in_297,
valid_in_298,valid_in_299,valid_in_300,valid_in_301,valid_in_302,valid_in_303,valid_in_304,valid_in_305,valid_in_306,
valid_in_307,valid_in_308,valid_in_309,valid_in_310,valid_in_311,valid_in_312,valid_in_313,valid_in_314,valid_in_315,
valid_in_316,valid_in_317,valid_in_318,valid_in_319,valid_in_320,valid_in_321,valid_in_322,valid_in_323,valid_in_324,
valid_in_325,valid_in_326,valid_in_327,valid_in_328,valid_in_329,valid_in_330,valid_in_331,valid_in_332,valid_in_333,
valid_in_334,valid_in_335,valid_in_336,valid_in_337,valid_in_338,valid_in_339,valid_in_340,valid_in_341,valid_in_342,
valid_in_343,valid_in_344,valid_in_345,valid_in_346,valid_in_347,valid_in_348,valid_in_349,valid_in_350,valid_in_351,
valid_in_352,valid_in_353,valid_in_354,valid_in_355,valid_in_356,valid_in_357,valid_in_358,valid_in_359,valid_in_360,
valid_in_361,valid_in_362,valid_in_363,valid_in_364,valid_in_365,valid_in_366,valid_in_367,valid_in_368,valid_in_369,
valid_in_370,valid_in_371,valid_in_372,valid_in_373,valid_in_374,valid_in_375,valid_in_376,valid_in_377,valid_in_378,
valid_in_379,valid_in_380,valid_in_381,valid_in_382,valid_in_383,valid_in_384,valid_in_385,valid_in_386,valid_in_387,
valid_in_388,valid_in_389,valid_in_390,valid_in_391,valid_in_392,valid_in_393,valid_in_394,valid_in_395,valid_in_396,
valid_in_397,valid_in_398,valid_in_399,valid_in_400,valid_in_401,valid_in_402,valid_in_403,valid_in_404,valid_in_405,
valid_in_406,valid_in_407,valid_in_408,valid_in_409,valid_in_410,valid_in_411,valid_in_412,valid_in_413,valid_in_414,
valid_in_415,valid_in_416,valid_in_417,valid_in_418,valid_in_419,valid_in_420,valid_in_421,valid_in_422,valid_in_423,
valid_in_424,valid_in_425,valid_in_426,valid_in_427,valid_in_428,valid_in_429,valid_in_430,valid_in_431,valid_in_432,
valid_in_433,valid_in_434,valid_in_435,valid_in_436,valid_in_437,valid_in_438,valid_in_439,valid_in_440,valid_in_441,
valid_in_442,valid_in_443,valid_in_444,valid_in_445,valid_in_446,valid_in_447,valid_in_448,valid_in_449,valid_in_450,
valid_in_451,valid_in_452,valid_in_453,valid_in_454,valid_in_455,valid_in_456,valid_in_457,valid_in_458,valid_in_459,
valid_in_460,valid_in_461,valid_in_462,valid_in_463,valid_in_464,valid_in_465,valid_in_466,valid_in_467,valid_in_468,
valid_in_469,valid_in_470,valid_in_471,valid_in_472,valid_in_473,valid_in_474,valid_in_475,valid_in_476,valid_in_477,
valid_in_478,valid_in_479,valid_in_480,valid_in_481,valid_in_482,valid_in_483,valid_in_484,valid_in_485,valid_in_486,
valid_in_487,valid_in_488,valid_in_489,valid_in_490,valid_in_491,valid_in_492,valid_in_493,valid_in_494,valid_in_495,
valid_in_496,valid_in_497,valid_in_498,valid_in_499,valid_in_500,valid_in_501,valid_in_502,valid_in_503,valid_in_504,
valid_in_505,valid_in_506,valid_in_507,valid_in_508,valid_in_509,valid_in_510,valid_in_511,valid_in_512,valid_in_513,
valid_in_514,valid_in_515,valid_in_516,valid_in_517,valid_in_518,valid_in_519,valid_in_520,valid_in_521,valid_in_522,
valid_in_523,valid_in_524,valid_in_525,valid_in_526,valid_in_527,valid_in_528,valid_in_529,valid_in_530,valid_in_531,
valid_in_532,valid_in_533,valid_in_534,valid_in_535,valid_in_536,valid_in_537,valid_in_538,valid_in_539,valid_in_540,
valid_in_541,valid_in_542,valid_in_543,valid_in_544,valid_in_545,valid_in_546,valid_in_547,valid_in_548,valid_in_549,
valid_in_550,valid_in_551,valid_in_552,valid_in_553,valid_in_554,valid_in_555,valid_in_556,valid_in_557,valid_in_558,
valid_in_559,valid_in_560,valid_in_561,valid_in_562,valid_in_563,valid_in_564,valid_in_565,valid_in_566,valid_in_567,
valid_in_568,valid_in_569,valid_in_570,valid_in_571,valid_in_572,valid_in_573,valid_in_574,valid_in_575,valid_in_576,
valid_in_577,valid_in_578,valid_in_579,valid_in_580,valid_in_581,valid_in_582,valid_in_583,valid_in_584,valid_in_585,
valid_in_586,valid_in_587,valid_in_588,valid_in_589,valid_in_590,valid_in_591,valid_in_592,valid_in_593,valid_in_594,
valid_in_595,valid_in_596,valid_in_597,valid_in_598,valid_in_599,valid_in_600,valid_in_601,valid_in_602,valid_in_603,
valid_in_604,valid_in_605,valid_in_606,valid_in_607,valid_in_608,valid_in_609,valid_in_610,valid_in_611,valid_in_612,
valid_in_613,valid_in_614,valid_in_615,valid_in_616,valid_in_617,valid_in_618,valid_in_619,valid_in_620,valid_in_621,
valid_in_622,valid_in_623,valid_in_624,valid_in_625,valid_in_626,valid_in_627,valid_in_628,valid_in_629,valid_in_630,
valid_in_631,valid_in_632,valid_in_633,valid_in_634,valid_in_635,valid_in_636,valid_in_637,valid_in_638,valid_in_639,
valid_in_640,valid_in_641,valid_in_642,valid_in_643,valid_in_644,valid_in_645,valid_in_646,valid_in_647,valid_in_648,
valid_in_649,valid_in_650,valid_in_651,valid_in_652,valid_in_653,valid_in_654,valid_in_655,valid_in_656,valid_in_657,
valid_in_658,valid_in_659,valid_in_660,valid_in_661,valid_in_662,valid_in_663,valid_in_664,valid_in_665,valid_in_666,
valid_in_667,valid_in_668,valid_in_669,valid_in_670,valid_in_671,valid_in_672,valid_in_673,valid_in_674,valid_in_675,
valid_in_676,valid_in_677,valid_in_678,valid_in_679,valid_in_680,valid_in_681,valid_in_682,valid_in_683,valid_in_684,
valid_in_685,valid_in_686,valid_in_687,valid_in_688,valid_in_689,valid_in_690,valid_in_691,valid_in_692,valid_in_693,
valid_in_694,valid_in_695,valid_in_696,valid_in_697,valid_in_698,valid_in_699,valid_in_700,valid_in_701,valid_in_702,
valid_in_703,valid_in_704,valid_in_705,valid_in_706,valid_in_707,valid_in_708,valid_in_709,valid_in_710,valid_in_711,
valid_in_712,valid_in_713,valid_in_714,valid_in_715,valid_in_716,valid_in_717,valid_in_718,valid_in_719,valid_in_720,
valid_in_721,valid_in_722,valid_in_723,valid_in_724,valid_in_725,valid_in_726,valid_in_727,valid_in_728,valid_in_729,
valid_in_730,valid_in_731,valid_in_732,valid_in_733,valid_in_734,valid_in_735,valid_in_736,valid_in_737,valid_in_738,
valid_in_739,valid_in_740,valid_in_741,valid_in_742,valid_in_743,valid_in_744,valid_in_745,valid_in_746,valid_in_747,
valid_in_748,valid_in_749,valid_in_750,valid_in_751,valid_in_752,valid_in_753,valid_in_754,valid_in_755,valid_in_756,
valid_in_757,valid_in_758,valid_in_759,valid_in_760,valid_in_761,valid_in_762,valid_in_763,valid_in_764,valid_in_765,
valid_in_766,valid_in_767,valid_in_768,valid_in_769,valid_in_770,valid_in_771,valid_in_772,valid_in_773,valid_in_774,
valid_in_775,valid_in_776,valid_in_777,valid_in_778,valid_in_779,valid_in_780,valid_in_781,valid_in_782,valid_in_783,
valid_in_784,valid_in_785,valid_in_786,valid_in_787,valid_in_788,valid_in_789,valid_in_790,valid_in_791,valid_in_792,
valid_in_793,valid_in_794,valid_in_795,valid_in_796,valid_in_797,valid_in_798,valid_in_799,valid_in_800,valid_in_801,
valid_in_802,valid_in_803,valid_in_804,valid_in_805,valid_in_806,valid_in_807,valid_in_808,valid_in_809,valid_in_810,
valid_in_811,valid_in_812,valid_in_813,valid_in_814,valid_in_815,valid_in_816,valid_in_817,valid_in_818,valid_in_819,
valid_in_820,valid_in_821,valid_in_822,valid_in_823,valid_in_824,valid_in_825,valid_in_826,valid_in_827,valid_in_828,
valid_in_829,valid_in_830,valid_in_831,valid_in_832,valid_in_833,valid_in_834,valid_in_835,valid_in_836,valid_in_837,
valid_in_838,valid_in_839,valid_in_840,valid_in_841,valid_in_842,valid_in_843,valid_in_844,valid_in_845,valid_in_846,
valid_in_847,valid_in_848,valid_in_849,valid_in_850,valid_in_851,valid_in_852,valid_in_853,valid_in_854,valid_in_855,
valid_in_856,valid_in_857,valid_in_858,valid_in_859,valid_in_860,valid_in_861,valid_in_862,valid_in_863,valid_in_864,
valid_in_865,valid_in_866,valid_in_867,valid_in_868,valid_in_869,valid_in_870,valid_in_871,valid_in_872,valid_in_873,
valid_in_874,valid_in_875,valid_in_876,valid_in_877,valid_in_878,valid_in_879,valid_in_880,valid_in_881,valid_in_882,
valid_in_883,valid_in_884,valid_in_885,valid_in_886,valid_in_887,valid_in_888,valid_in_889,valid_in_890,valid_in_891,
valid_in_892,valid_in_893,valid_in_894,valid_in_895,valid_in_896,valid_in_897,valid_in_898,valid_in_899,valid_in_900,
valid_in_901,valid_in_902,valid_in_903,valid_in_904,valid_in_905,valid_in_906,valid_in_907,valid_in_908,valid_in_909,
valid_in_910,valid_in_911,valid_in_912,valid_in_913,valid_in_914,valid_in_915,valid_in_916,valid_in_917,valid_in_918,
valid_in_919,valid_in_920,valid_in_921,valid_in_922,valid_in_923,valid_in_924,valid_in_925,valid_in_926,valid_in_927,
valid_in_928,valid_in_929,valid_in_930,valid_in_931,valid_in_932,valid_in_933,valid_in_934,valid_in_935,valid_in_936,
valid_in_937,valid_in_938,valid_in_939,valid_in_940,valid_in_941,valid_in_942,valid_in_943,valid_in_944,valid_in_945,
valid_in_946,valid_in_947,valid_in_948,valid_in_949,valid_in_950,valid_in_951,valid_in_952,valid_in_953,valid_in_954,
valid_in_955,valid_in_956,valid_in_957,valid_in_958,valid_in_959,valid_in_960,valid_in_961,valid_in_962,valid_in_963,
valid_in_964,valid_in_965,valid_in_966,valid_in_967,valid_in_968,valid_in_969,valid_in_970,valid_in_971,valid_in_972,
valid_in_973,valid_in_974,valid_in_975,valid_in_976,valid_in_977,valid_in_978,valid_in_979,valid_in_980,valid_in_981,
valid_in_982,valid_in_983,valid_in_984,valid_in_985,valid_in_986,valid_in_987,valid_in_988,valid_in_989,valid_in_990,
valid_in_991,valid_in_992,valid_in_993,valid_in_994,valid_in_995,valid_in_996,valid_in_997,valid_in_998,valid_in_999,
valid_in_1000,valid_in_1001,valid_in_1002,valid_in_1003,valid_in_1004,valid_in_1005,valid_in_1006,valid_in_1007,valid_in_1008,
valid_in_1009,valid_in_1010,valid_in_1011,valid_in_1012,valid_in_1013,valid_in_1014,valid_in_1015,valid_in_1016,valid_in_1017,
valid_in_1018,valid_in_1019,valid_in_1020,valid_in_1021,valid_in_1022,valid_in_1023,valid_in_1024,
    	      
    	input [DATA_WIDTH-1:0] pxl_in_1,pxl_in_2,pxl_in_3,pxl_in_4,pxl_in_5,pxl_in_6,pxl_in_7,pxl_in_8,pxl_in_9,
pxl_in_10,pxl_in_11,pxl_in_12,pxl_in_13,pxl_in_14,pxl_in_15,pxl_in_16,pxl_in_17,pxl_in_18,
pxl_in_19,pxl_in_20,pxl_in_21,pxl_in_22,pxl_in_23,pxl_in_24,pxl_in_25,pxl_in_26,pxl_in_27,
pxl_in_28,pxl_in_29,pxl_in_30,pxl_in_31,pxl_in_32,pxl_in_33,pxl_in_34,pxl_in_35,pxl_in_36,
pxl_in_37,pxl_in_38,pxl_in_39,pxl_in_40,pxl_in_41,pxl_in_42,pxl_in_43,pxl_in_44,pxl_in_45,
pxl_in_46,pxl_in_47,pxl_in_48,pxl_in_49,pxl_in_50,pxl_in_51,pxl_in_52,pxl_in_53,pxl_in_54,
pxl_in_55,pxl_in_56,pxl_in_57,pxl_in_58,pxl_in_59,pxl_in_60,pxl_in_61,pxl_in_62,pxl_in_63,
pxl_in_64,pxl_in_65,pxl_in_66,pxl_in_67,pxl_in_68,pxl_in_69,pxl_in_70,pxl_in_71,pxl_in_72,
pxl_in_73,pxl_in_74,pxl_in_75,pxl_in_76,pxl_in_77,pxl_in_78,pxl_in_79,pxl_in_80,pxl_in_81,
pxl_in_82,pxl_in_83,pxl_in_84,pxl_in_85,pxl_in_86,pxl_in_87,pxl_in_88,pxl_in_89,pxl_in_90,
pxl_in_91,pxl_in_92,pxl_in_93,pxl_in_94,pxl_in_95,pxl_in_96,pxl_in_97,pxl_in_98,pxl_in_99,
pxl_in_100,pxl_in_101,pxl_in_102,pxl_in_103,pxl_in_104,pxl_in_105,pxl_in_106,pxl_in_107,pxl_in_108,
pxl_in_109,pxl_in_110,pxl_in_111,pxl_in_112,pxl_in_113,pxl_in_114,pxl_in_115,pxl_in_116,pxl_in_117,
pxl_in_118,pxl_in_119,pxl_in_120,pxl_in_121,pxl_in_122,pxl_in_123,pxl_in_124,pxl_in_125,pxl_in_126,
pxl_in_127,pxl_in_128,pxl_in_129,pxl_in_130,pxl_in_131,pxl_in_132,pxl_in_133,pxl_in_134,pxl_in_135,
pxl_in_136,pxl_in_137,pxl_in_138,pxl_in_139,pxl_in_140,pxl_in_141,pxl_in_142,pxl_in_143,pxl_in_144,
pxl_in_145,pxl_in_146,pxl_in_147,pxl_in_148,pxl_in_149,pxl_in_150,pxl_in_151,pxl_in_152,pxl_in_153,
pxl_in_154,pxl_in_155,pxl_in_156,pxl_in_157,pxl_in_158,pxl_in_159,pxl_in_160,pxl_in_161,pxl_in_162,
pxl_in_163,pxl_in_164,pxl_in_165,pxl_in_166,pxl_in_167,pxl_in_168,pxl_in_169,pxl_in_170,pxl_in_171,
pxl_in_172,pxl_in_173,pxl_in_174,pxl_in_175,pxl_in_176,pxl_in_177,pxl_in_178,pxl_in_179,pxl_in_180,
pxl_in_181,pxl_in_182,pxl_in_183,pxl_in_184,pxl_in_185,pxl_in_186,pxl_in_187,pxl_in_188,pxl_in_189,
pxl_in_190,pxl_in_191,pxl_in_192,pxl_in_193,pxl_in_194,pxl_in_195,pxl_in_196,pxl_in_197,pxl_in_198,
pxl_in_199,pxl_in_200,pxl_in_201,pxl_in_202,pxl_in_203,pxl_in_204,pxl_in_205,pxl_in_206,pxl_in_207,
pxl_in_208,pxl_in_209,pxl_in_210,pxl_in_211,pxl_in_212,pxl_in_213,pxl_in_214,pxl_in_215,pxl_in_216,
pxl_in_217,pxl_in_218,pxl_in_219,pxl_in_220,pxl_in_221,pxl_in_222,pxl_in_223,pxl_in_224,pxl_in_225,
pxl_in_226,pxl_in_227,pxl_in_228,pxl_in_229,pxl_in_230,pxl_in_231,pxl_in_232,pxl_in_233,pxl_in_234,
pxl_in_235,pxl_in_236,pxl_in_237,pxl_in_238,pxl_in_239,pxl_in_240,pxl_in_241,pxl_in_242,pxl_in_243,
pxl_in_244,pxl_in_245,pxl_in_246,pxl_in_247,pxl_in_248,pxl_in_249,pxl_in_250,pxl_in_251,pxl_in_252,
pxl_in_253,pxl_in_254,pxl_in_255,pxl_in_256,pxl_in_257,pxl_in_258,pxl_in_259,pxl_in_260,pxl_in_261,
pxl_in_262,pxl_in_263,pxl_in_264,pxl_in_265,pxl_in_266,pxl_in_267,pxl_in_268,pxl_in_269,pxl_in_270,
pxl_in_271,pxl_in_272,pxl_in_273,pxl_in_274,pxl_in_275,pxl_in_276,pxl_in_277,pxl_in_278,pxl_in_279,
pxl_in_280,pxl_in_281,pxl_in_282,pxl_in_283,pxl_in_284,pxl_in_285,pxl_in_286,pxl_in_287,pxl_in_288,
pxl_in_289,pxl_in_290,pxl_in_291,pxl_in_292,pxl_in_293,pxl_in_294,pxl_in_295,pxl_in_296,pxl_in_297,
pxl_in_298,pxl_in_299,pxl_in_300,pxl_in_301,pxl_in_302,pxl_in_303,pxl_in_304,pxl_in_305,pxl_in_306,
pxl_in_307,pxl_in_308,pxl_in_309,pxl_in_310,pxl_in_311,pxl_in_312,pxl_in_313,pxl_in_314,pxl_in_315,
pxl_in_316,pxl_in_317,pxl_in_318,pxl_in_319,pxl_in_320,pxl_in_321,pxl_in_322,pxl_in_323,pxl_in_324,
pxl_in_325,pxl_in_326,pxl_in_327,pxl_in_328,pxl_in_329,pxl_in_330,pxl_in_331,pxl_in_332,pxl_in_333,
pxl_in_334,pxl_in_335,pxl_in_336,pxl_in_337,pxl_in_338,pxl_in_339,pxl_in_340,pxl_in_341,pxl_in_342,
pxl_in_343,pxl_in_344,pxl_in_345,pxl_in_346,pxl_in_347,pxl_in_348,pxl_in_349,pxl_in_350,pxl_in_351,
pxl_in_352,pxl_in_353,pxl_in_354,pxl_in_355,pxl_in_356,pxl_in_357,pxl_in_358,pxl_in_359,pxl_in_360,
pxl_in_361,pxl_in_362,pxl_in_363,pxl_in_364,pxl_in_365,pxl_in_366,pxl_in_367,pxl_in_368,pxl_in_369,
pxl_in_370,pxl_in_371,pxl_in_372,pxl_in_373,pxl_in_374,pxl_in_375,pxl_in_376,pxl_in_377,pxl_in_378,
pxl_in_379,pxl_in_380,pxl_in_381,pxl_in_382,pxl_in_383,pxl_in_384,pxl_in_385,pxl_in_386,pxl_in_387,
pxl_in_388,pxl_in_389,pxl_in_390,pxl_in_391,pxl_in_392,pxl_in_393,pxl_in_394,pxl_in_395,pxl_in_396,
pxl_in_397,pxl_in_398,pxl_in_399,pxl_in_400,pxl_in_401,pxl_in_402,pxl_in_403,pxl_in_404,pxl_in_405,
pxl_in_406,pxl_in_407,pxl_in_408,pxl_in_409,pxl_in_410,pxl_in_411,pxl_in_412,pxl_in_413,pxl_in_414,
pxl_in_415,pxl_in_416,pxl_in_417,pxl_in_418,pxl_in_419,pxl_in_420,pxl_in_421,pxl_in_422,pxl_in_423,
pxl_in_424,pxl_in_425,pxl_in_426,pxl_in_427,pxl_in_428,pxl_in_429,pxl_in_430,pxl_in_431,pxl_in_432,
pxl_in_433,pxl_in_434,pxl_in_435,pxl_in_436,pxl_in_437,pxl_in_438,pxl_in_439,pxl_in_440,pxl_in_441,
pxl_in_442,pxl_in_443,pxl_in_444,pxl_in_445,pxl_in_446,pxl_in_447,pxl_in_448,pxl_in_449,pxl_in_450,
pxl_in_451,pxl_in_452,pxl_in_453,pxl_in_454,pxl_in_455,pxl_in_456,pxl_in_457,pxl_in_458,pxl_in_459,
pxl_in_460,pxl_in_461,pxl_in_462,pxl_in_463,pxl_in_464,pxl_in_465,pxl_in_466,pxl_in_467,pxl_in_468,
pxl_in_469,pxl_in_470,pxl_in_471,pxl_in_472,pxl_in_473,pxl_in_474,pxl_in_475,pxl_in_476,pxl_in_477,
pxl_in_478,pxl_in_479,pxl_in_480,pxl_in_481,pxl_in_482,pxl_in_483,pxl_in_484,pxl_in_485,pxl_in_486,
pxl_in_487,pxl_in_488,pxl_in_489,pxl_in_490,pxl_in_491,pxl_in_492,pxl_in_493,pxl_in_494,pxl_in_495,
pxl_in_496,pxl_in_497,pxl_in_498,pxl_in_499,pxl_in_500,pxl_in_501,pxl_in_502,pxl_in_503,pxl_in_504,
pxl_in_505,pxl_in_506,pxl_in_507,pxl_in_508,pxl_in_509,pxl_in_510,pxl_in_511,pxl_in_512,pxl_in_513,
pxl_in_514,pxl_in_515,pxl_in_516,pxl_in_517,pxl_in_518,pxl_in_519,pxl_in_520,pxl_in_521,pxl_in_522,
pxl_in_523,pxl_in_524,pxl_in_525,pxl_in_526,pxl_in_527,pxl_in_528,pxl_in_529,pxl_in_530,pxl_in_531,
pxl_in_532,pxl_in_533,pxl_in_534,pxl_in_535,pxl_in_536,pxl_in_537,pxl_in_538,pxl_in_539,pxl_in_540,
pxl_in_541,pxl_in_542,pxl_in_543,pxl_in_544,pxl_in_545,pxl_in_546,pxl_in_547,pxl_in_548,pxl_in_549,
pxl_in_550,pxl_in_551,pxl_in_552,pxl_in_553,pxl_in_554,pxl_in_555,pxl_in_556,pxl_in_557,pxl_in_558,
pxl_in_559,pxl_in_560,pxl_in_561,pxl_in_562,pxl_in_563,pxl_in_564,pxl_in_565,pxl_in_566,pxl_in_567,
pxl_in_568,pxl_in_569,pxl_in_570,pxl_in_571,pxl_in_572,pxl_in_573,pxl_in_574,pxl_in_575,pxl_in_576,
pxl_in_577,pxl_in_578,pxl_in_579,pxl_in_580,pxl_in_581,pxl_in_582,pxl_in_583,pxl_in_584,pxl_in_585,
pxl_in_586,pxl_in_587,pxl_in_588,pxl_in_589,pxl_in_590,pxl_in_591,pxl_in_592,pxl_in_593,pxl_in_594,
pxl_in_595,pxl_in_596,pxl_in_597,pxl_in_598,pxl_in_599,pxl_in_600,pxl_in_601,pxl_in_602,pxl_in_603,
pxl_in_604,pxl_in_605,pxl_in_606,pxl_in_607,pxl_in_608,pxl_in_609,pxl_in_610,pxl_in_611,pxl_in_612,
pxl_in_613,pxl_in_614,pxl_in_615,pxl_in_616,pxl_in_617,pxl_in_618,pxl_in_619,pxl_in_620,pxl_in_621,
pxl_in_622,pxl_in_623,pxl_in_624,pxl_in_625,pxl_in_626,pxl_in_627,pxl_in_628,pxl_in_629,pxl_in_630,
pxl_in_631,pxl_in_632,pxl_in_633,pxl_in_634,pxl_in_635,pxl_in_636,pxl_in_637,pxl_in_638,pxl_in_639,
pxl_in_640,pxl_in_641,pxl_in_642,pxl_in_643,pxl_in_644,pxl_in_645,pxl_in_646,pxl_in_647,pxl_in_648,
pxl_in_649,pxl_in_650,pxl_in_651,pxl_in_652,pxl_in_653,pxl_in_654,pxl_in_655,pxl_in_656,pxl_in_657,
pxl_in_658,pxl_in_659,pxl_in_660,pxl_in_661,pxl_in_662,pxl_in_663,pxl_in_664,pxl_in_665,pxl_in_666,
pxl_in_667,pxl_in_668,pxl_in_669,pxl_in_670,pxl_in_671,pxl_in_672,pxl_in_673,pxl_in_674,pxl_in_675,
pxl_in_676,pxl_in_677,pxl_in_678,pxl_in_679,pxl_in_680,pxl_in_681,pxl_in_682,pxl_in_683,pxl_in_684,
pxl_in_685,pxl_in_686,pxl_in_687,pxl_in_688,pxl_in_689,pxl_in_690,pxl_in_691,pxl_in_692,pxl_in_693,
pxl_in_694,pxl_in_695,pxl_in_696,pxl_in_697,pxl_in_698,pxl_in_699,pxl_in_700,pxl_in_701,pxl_in_702,
pxl_in_703,pxl_in_704,pxl_in_705,pxl_in_706,pxl_in_707,pxl_in_708,pxl_in_709,pxl_in_710,pxl_in_711,
pxl_in_712,pxl_in_713,pxl_in_714,pxl_in_715,pxl_in_716,pxl_in_717,pxl_in_718,pxl_in_719,pxl_in_720,
pxl_in_721,pxl_in_722,pxl_in_723,pxl_in_724,pxl_in_725,pxl_in_726,pxl_in_727,pxl_in_728,pxl_in_729,
pxl_in_730,pxl_in_731,pxl_in_732,pxl_in_733,pxl_in_734,pxl_in_735,pxl_in_736,pxl_in_737,pxl_in_738,
pxl_in_739,pxl_in_740,pxl_in_741,pxl_in_742,pxl_in_743,pxl_in_744,pxl_in_745,pxl_in_746,pxl_in_747,
pxl_in_748,pxl_in_749,pxl_in_750,pxl_in_751,pxl_in_752,pxl_in_753,pxl_in_754,pxl_in_755,pxl_in_756,
pxl_in_757,pxl_in_758,pxl_in_759,pxl_in_760,pxl_in_761,pxl_in_762,pxl_in_763,pxl_in_764,pxl_in_765,
pxl_in_766,pxl_in_767,pxl_in_768,pxl_in_769,pxl_in_770,pxl_in_771,pxl_in_772,pxl_in_773,pxl_in_774,
pxl_in_775,pxl_in_776,pxl_in_777,pxl_in_778,pxl_in_779,pxl_in_780,pxl_in_781,pxl_in_782,pxl_in_783,
pxl_in_784,pxl_in_785,pxl_in_786,pxl_in_787,pxl_in_788,pxl_in_789,pxl_in_790,pxl_in_791,pxl_in_792,
pxl_in_793,pxl_in_794,pxl_in_795,pxl_in_796,pxl_in_797,pxl_in_798,pxl_in_799,pxl_in_800,pxl_in_801,
pxl_in_802,pxl_in_803,pxl_in_804,pxl_in_805,pxl_in_806,pxl_in_807,pxl_in_808,pxl_in_809,pxl_in_810,
pxl_in_811,pxl_in_812,pxl_in_813,pxl_in_814,pxl_in_815,pxl_in_816,pxl_in_817,pxl_in_818,pxl_in_819,
pxl_in_820,pxl_in_821,pxl_in_822,pxl_in_823,pxl_in_824,pxl_in_825,pxl_in_826,pxl_in_827,pxl_in_828,
pxl_in_829,pxl_in_830,pxl_in_831,pxl_in_832,pxl_in_833,pxl_in_834,pxl_in_835,pxl_in_836,pxl_in_837,
pxl_in_838,pxl_in_839,pxl_in_840,pxl_in_841,pxl_in_842,pxl_in_843,pxl_in_844,pxl_in_845,pxl_in_846,
pxl_in_847,pxl_in_848,pxl_in_849,pxl_in_850,pxl_in_851,pxl_in_852,pxl_in_853,pxl_in_854,pxl_in_855,
pxl_in_856,pxl_in_857,pxl_in_858,pxl_in_859,pxl_in_860,pxl_in_861,pxl_in_862,pxl_in_863,pxl_in_864,
pxl_in_865,pxl_in_866,pxl_in_867,pxl_in_868,pxl_in_869,pxl_in_870,pxl_in_871,pxl_in_872,pxl_in_873,
pxl_in_874,pxl_in_875,pxl_in_876,pxl_in_877,pxl_in_878,pxl_in_879,pxl_in_880,pxl_in_881,pxl_in_882,
pxl_in_883,pxl_in_884,pxl_in_885,pxl_in_886,pxl_in_887,pxl_in_888,pxl_in_889,pxl_in_890,pxl_in_891,
pxl_in_892,pxl_in_893,pxl_in_894,pxl_in_895,pxl_in_896,pxl_in_897,pxl_in_898,pxl_in_899,pxl_in_900,
pxl_in_901,pxl_in_902,pxl_in_903,pxl_in_904,pxl_in_905,pxl_in_906,pxl_in_907,pxl_in_908,pxl_in_909,
pxl_in_910,pxl_in_911,pxl_in_912,pxl_in_913,pxl_in_914,pxl_in_915,pxl_in_916,pxl_in_917,pxl_in_918,
pxl_in_919,pxl_in_920,pxl_in_921,pxl_in_922,pxl_in_923,pxl_in_924,pxl_in_925,pxl_in_926,pxl_in_927,
pxl_in_928,pxl_in_929,pxl_in_930,pxl_in_931,pxl_in_932,pxl_in_933,pxl_in_934,pxl_in_935,pxl_in_936,
pxl_in_937,pxl_in_938,pxl_in_939,pxl_in_940,pxl_in_941,pxl_in_942,pxl_in_943,pxl_in_944,pxl_in_945,
pxl_in_946,pxl_in_947,pxl_in_948,pxl_in_949,pxl_in_950,pxl_in_951,pxl_in_952,pxl_in_953,pxl_in_954,
pxl_in_955,pxl_in_956,pxl_in_957,pxl_in_958,pxl_in_959,pxl_in_960,pxl_in_961,pxl_in_962,pxl_in_963,
pxl_in_964,pxl_in_965,pxl_in_966,pxl_in_967,pxl_in_968,pxl_in_969,pxl_in_970,pxl_in_971,pxl_in_972,
pxl_in_973,pxl_in_974,pxl_in_975,pxl_in_976,pxl_in_977,pxl_in_978,pxl_in_979,pxl_in_980,pxl_in_981,
pxl_in_982,pxl_in_983,pxl_in_984,pxl_in_985,pxl_in_986,pxl_in_987,pxl_in_988,pxl_in_989,pxl_in_990,
pxl_in_991,pxl_in_992,pxl_in_993,pxl_in_994,pxl_in_995,pxl_in_996,pxl_in_997,pxl_in_998,pxl_in_999,
pxl_in_1000,pxl_in_1001,pxl_in_1002,pxl_in_1003,pxl_in_1004,pxl_in_1005,pxl_in_1006,pxl_in_1007,pxl_in_1008,
pxl_in_1009,pxl_in_1010,pxl_in_1011,pxl_in_1012,pxl_in_1013,pxl_in_1014,pxl_in_1015,pxl_in_1016,pxl_in_1017,
pxl_in_1018,pxl_in_1019,pxl_in_1020,pxl_in_1021,pxl_in_1022,pxl_in_1023,pxl_in_1024,
  	     	
    	output [DATA_WIDTH-1:0] pxl_out_1 , pxl_out_2 , pxl_out_3 , pxl_out_4 , pxl_out_5 , pxl_out_6 , pxl_out_7 , pxl_out_8 , pxl_out_9 , pxl_out_10,
                        pxl_out_11, pxl_out_12, pxl_out_13, pxl_out_14, pxl_out_15, pxl_out_16, pxl_out_17, pxl_out_18, pxl_out_19, pxl_out_20,
	                      pxl_out_21, pxl_out_22, pxl_out_23, pxl_out_24, pxl_out_25, pxl_out_26, pxl_out_27, pxl_out_28, pxl_out_29, pxl_out_30,
                        pxl_out_31, pxl_out_32,
	                                 
	               output valid_out_1 , valid_out_2 , valid_out_3 , valid_out_4 , valid_out_5 , valid_out_6 , valid_out_7 , valid_out_8 , valid_out_9 , valid_out_10,
                        valid_out_11, valid_out_12, valid_out_13, valid_out_14, valid_out_15, valid_out_16, valid_out_17, valid_out_18, valid_out_19, valid_out_20,
	                      valid_out_21, valid_out_22, valid_out_23, valid_out_24, valid_out_25, valid_out_26, valid_out_27, valid_out_28, valid_out_29, valid_out_30,
                        valid_out_31, valid_out_32
	 );
	 
add_32layers#(D, DATA_WIDTH) x1(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_1), .pxl_in_1(pxl_in_1), .valid_in_2(valid_in_2), .pxl_in_2(pxl_in_2), .valid_in_3(valid_in_3), .pxl_in_3(pxl_in_3), .valid_in_4(valid_in_4), .pxl_in_4(pxl_in_4), .valid_in_5(valid_in_5), .pxl_in_5(pxl_in_5), .valid_in_6(valid_in_6), .pxl_in_6(pxl_in_6), .valid_in_7(valid_in_7), .pxl_in_7(pxl_in_7), .valid_in_8(valid_in_8), .pxl_in_8(pxl_in_8), .valid_in_9(valid_in_9), .pxl_in_9(pxl_in_9), .valid_in_10(valid_in_10), .pxl_in_10(pxl_in_10), .valid_in_11(valid_in_11), .pxl_in_11(pxl_in_11), .valid_in_12(valid_in_12), .pxl_in_12(pxl_in_12), .valid_in_13(valid_in_13), .pxl_in_13(pxl_in_13), .valid_in_14(valid_in_14), .pxl_in_14(pxl_in_14), .valid_in_15(valid_in_15), .pxl_in_15(pxl_in_15), .valid_in_16(valid_in_16), .pxl_in_16(pxl_in_16), .valid_in_17(valid_in_17), .pxl_in_17(pxl_in_17), .valid_in_18(valid_in_18), .pxl_in_18(pxl_in_18), .valid_in_19(valid_in_19), .pxl_in_19(pxl_in_19), .valid_in_20(valid_in_20), .pxl_in_20(pxl_in_20), .valid_in_21(valid_in_21), .pxl_in_21(pxl_in_21), .valid_in_22(valid_in_22), .pxl_in_22(pxl_in_22), .valid_in_23(valid_in_23), .pxl_in_23(pxl_in_23), .valid_in_24(valid_in_24), .pxl_in_24(pxl_in_24), .valid_in_25(valid_in_25), .pxl_in_25(pxl_in_25), .valid_in_26(valid_in_26), .pxl_in_26(pxl_in_26), .valid_in_27(valid_in_27), .pxl_in_27(pxl_in_27), .valid_in_28(valid_in_28), .pxl_in_28(pxl_in_28), .valid_in_29(valid_in_29), .pxl_in_29(pxl_in_29), .valid_in_30(valid_in_30), .pxl_in_30(pxl_in_30), .valid_in_31(valid_in_31), .pxl_in_31(pxl_in_31), .valid_in_32(valid_in_32), .pxl_in_32(pxl_in_32), .pxl_out(pxl_out_1), .valid_out(valid_out_1) );

add_32layers#(D, DATA_WIDTH) x2(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_33), .pxl_in_1(pxl_in_33), .valid_in_2(valid_in_34), .pxl_in_2(pxl_in_34), .valid_in_3(valid_in_35), .pxl_in_3(pxl_in_35), .valid_in_4(valid_in_36), .pxl_in_4(pxl_in_36), .valid_in_5(valid_in_37), .pxl_in_5(pxl_in_37), .valid_in_6(valid_in_38), .pxl_in_6(pxl_in_38), .valid_in_7(valid_in_39), .pxl_in_7(pxl_in_39), .valid_in_8(valid_in_40), .pxl_in_8(pxl_in_40), .valid_in_9(valid_in_41), .pxl_in_9(pxl_in_41), .valid_in_10(valid_in_42), .pxl_in_10(pxl_in_42), .valid_in_11(valid_in_43), .pxl_in_11(pxl_in_43), .valid_in_12(valid_in_44), .pxl_in_12(pxl_in_44), .valid_in_13(valid_in_45), .pxl_in_13(pxl_in_45), .valid_in_14(valid_in_46), .pxl_in_14(pxl_in_46), .valid_in_15(valid_in_47), .pxl_in_15(pxl_in_47), .valid_in_16(valid_in_48), .pxl_in_16(pxl_in_48), .valid_in_17(valid_in_49), .pxl_in_17(pxl_in_49), .valid_in_18(valid_in_50), .pxl_in_18(pxl_in_50), .valid_in_19(valid_in_51), .pxl_in_19(pxl_in_51), .valid_in_20(valid_in_52), .pxl_in_20(pxl_in_52), .valid_in_21(valid_in_53), .pxl_in_21(pxl_in_53), .valid_in_22(valid_in_54), .pxl_in_22(pxl_in_54), .valid_in_23(valid_in_55), .pxl_in_23(pxl_in_55), .valid_in_24(valid_in_56), .pxl_in_24(pxl_in_56), .valid_in_25(valid_in_57), .pxl_in_25(pxl_in_57), .valid_in_26(valid_in_58), .pxl_in_26(pxl_in_58), .valid_in_27(valid_in_59), .pxl_in_27(pxl_in_59), .valid_in_28(valid_in_60), .pxl_in_28(pxl_in_60), .valid_in_29(valid_in_61), .pxl_in_29(pxl_in_61), .valid_in_30(valid_in_62), .pxl_in_30(pxl_in_62), .valid_in_31(valid_in_63), .pxl_in_31(pxl_in_63), .valid_in_32(valid_in_64), .pxl_in_32(pxl_in_64), .pxl_out(pxl_out_2), .valid_out(valid_out_2) );

add_32layers#(D, DATA_WIDTH) x3(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_65), .pxl_in_1(pxl_in_65), .valid_in_2(valid_in_66), .pxl_in_2(pxl_in_66), .valid_in_3(valid_in_67), .pxl_in_3(pxl_in_67), .valid_in_4(valid_in_68), .pxl_in_4(pxl_in_68), .valid_in_5(valid_in_69), .pxl_in_5(pxl_in_69), .valid_in_6(valid_in_70), .pxl_in_6(pxl_in_70), .valid_in_7(valid_in_71), .pxl_in_7(pxl_in_71), .valid_in_8(valid_in_72), .pxl_in_8(pxl_in_72), .valid_in_9(valid_in_73), .pxl_in_9(pxl_in_73), .valid_in_10(valid_in_74), .pxl_in_10(pxl_in_74), .valid_in_11(valid_in_75), .pxl_in_11(pxl_in_75), .valid_in_12(valid_in_76), .pxl_in_12(pxl_in_76), .valid_in_13(valid_in_77), .pxl_in_13(pxl_in_77), .valid_in_14(valid_in_78), .pxl_in_14(pxl_in_78), .valid_in_15(valid_in_79), .pxl_in_15(pxl_in_79), .valid_in_16(valid_in_80), .pxl_in_16(pxl_in_80), .valid_in_17(valid_in_81), .pxl_in_17(pxl_in_81), .valid_in_18(valid_in_82), .pxl_in_18(pxl_in_82), .valid_in_19(valid_in_83), .pxl_in_19(pxl_in_83), .valid_in_20(valid_in_84), .pxl_in_20(pxl_in_84), .valid_in_21(valid_in_85), .pxl_in_21(pxl_in_85), .valid_in_22(valid_in_86), .pxl_in_22(pxl_in_86), .valid_in_23(valid_in_87), .pxl_in_23(pxl_in_87), .valid_in_24(valid_in_88), .pxl_in_24(pxl_in_88), .valid_in_25(valid_in_89), .pxl_in_25(pxl_in_89), .valid_in_26(valid_in_90), .pxl_in_26(pxl_in_90), .valid_in_27(valid_in_91), .pxl_in_27(pxl_in_91), .valid_in_28(valid_in_92), .pxl_in_28(pxl_in_92), .valid_in_29(valid_in_93), .pxl_in_29(pxl_in_93), .valid_in_30(valid_in_94), .pxl_in_30(pxl_in_94), .valid_in_31(valid_in_95), .pxl_in_31(pxl_in_95), .valid_in_32(valid_in_96), .pxl_in_32(pxl_in_96), .pxl_out(pxl_out_3), .valid_out(valid_out_3) );

add_32layers#(D, DATA_WIDTH) x4(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_97), .pxl_in_1(pxl_in_97), .valid_in_2(valid_in_98), .pxl_in_2(pxl_in_98), .valid_in_3(valid_in_99), .pxl_in_3(pxl_in_99), .valid_in_4(valid_in_100), .pxl_in_4(pxl_in_100), .valid_in_5(valid_in_101), .pxl_in_5(pxl_in_101), .valid_in_6(valid_in_102), .pxl_in_6(pxl_in_102), .valid_in_7(valid_in_103), .pxl_in_7(pxl_in_103), .valid_in_8(valid_in_104), .pxl_in_8(pxl_in_104), .valid_in_9(valid_in_105), .pxl_in_9(pxl_in_105), .valid_in_10(valid_in_106), .pxl_in_10(pxl_in_106), .valid_in_11(valid_in_107), .pxl_in_11(pxl_in_107), .valid_in_12(valid_in_108), .pxl_in_12(pxl_in_108), .valid_in_13(valid_in_109), .pxl_in_13(pxl_in_109), .valid_in_14(valid_in_110), .pxl_in_14(pxl_in_110), .valid_in_15(valid_in_111), .pxl_in_15(pxl_in_111), .valid_in_16(valid_in_112), .pxl_in_16(pxl_in_112), .valid_in_17(valid_in_113), .pxl_in_17(pxl_in_113), .valid_in_18(valid_in_114), .pxl_in_18(pxl_in_114), .valid_in_19(valid_in_115), .pxl_in_19(pxl_in_115), .valid_in_20(valid_in_116), .pxl_in_20(pxl_in_116), .valid_in_21(valid_in_117), .pxl_in_21(pxl_in_117), .valid_in_22(valid_in_118), .pxl_in_22(pxl_in_118), .valid_in_23(valid_in_119), .pxl_in_23(pxl_in_119), .valid_in_24(valid_in_120), .pxl_in_24(pxl_in_120), .valid_in_25(valid_in_121), .pxl_in_25(pxl_in_121), .valid_in_26(valid_in_122), .pxl_in_26(pxl_in_122), .valid_in_27(valid_in_123), .pxl_in_27(pxl_in_123), .valid_in_28(valid_in_124), .pxl_in_28(pxl_in_124), .valid_in_29(valid_in_125), .pxl_in_29(pxl_in_125), .valid_in_30(valid_in_126), .pxl_in_30(pxl_in_126), .valid_in_31(valid_in_127), .pxl_in_31(pxl_in_127), .valid_in_32(valid_in_128), .pxl_in_32(pxl_in_128), .pxl_out(pxl_out_4), .valid_out(valid_out_4) );

add_32layers#(D, DATA_WIDTH) x5(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_129), .pxl_in_1(pxl_in_129), .valid_in_2(valid_in_130), .pxl_in_2(pxl_in_130), .valid_in_3(valid_in_131), .pxl_in_3(pxl_in_131), .valid_in_4(valid_in_132), .pxl_in_4(pxl_in_132), .valid_in_5(valid_in_133), .pxl_in_5(pxl_in_133), .valid_in_6(valid_in_134), .pxl_in_6(pxl_in_134), .valid_in_7(valid_in_135), .pxl_in_7(pxl_in_135), .valid_in_8(valid_in_136), .pxl_in_8(pxl_in_136), .valid_in_9(valid_in_137), .pxl_in_9(pxl_in_137), .valid_in_10(valid_in_138), .pxl_in_10(pxl_in_138), .valid_in_11(valid_in_139), .pxl_in_11(pxl_in_139), .valid_in_12(valid_in_140), .pxl_in_12(pxl_in_140), .valid_in_13(valid_in_141), .pxl_in_13(pxl_in_141), .valid_in_14(valid_in_142), .pxl_in_14(pxl_in_142), .valid_in_15(valid_in_143), .pxl_in_15(pxl_in_143), .valid_in_16(valid_in_144), .pxl_in_16(pxl_in_144), .valid_in_17(valid_in_145), .pxl_in_17(pxl_in_145), .valid_in_18(valid_in_146), .pxl_in_18(pxl_in_146), .valid_in_19(valid_in_147), .pxl_in_19(pxl_in_147), .valid_in_20(valid_in_148), .pxl_in_20(pxl_in_148), .valid_in_21(valid_in_149), .pxl_in_21(pxl_in_149), .valid_in_22(valid_in_150), .pxl_in_22(pxl_in_150), .valid_in_23(valid_in_151), .pxl_in_23(pxl_in_151), .valid_in_24(valid_in_152), .pxl_in_24(pxl_in_152), .valid_in_25(valid_in_153), .pxl_in_25(pxl_in_153), .valid_in_26(valid_in_154), .pxl_in_26(pxl_in_154), .valid_in_27(valid_in_155), .pxl_in_27(pxl_in_155), .valid_in_28(valid_in_156), .pxl_in_28(pxl_in_156), .valid_in_29(valid_in_157), .pxl_in_29(pxl_in_157), .valid_in_30(valid_in_158), .pxl_in_30(pxl_in_158), .valid_in_31(valid_in_159), .pxl_in_31(pxl_in_159), .valid_in_32(valid_in_160), .pxl_in_32(pxl_in_160), .pxl_out(pxl_out_5), .valid_out(valid_out_5) );

add_32layers#(D, DATA_WIDTH) x6(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_161), .pxl_in_1(pxl_in_161), .valid_in_2(valid_in_162), .pxl_in_2(pxl_in_162), .valid_in_3(valid_in_163), .pxl_in_3(pxl_in_163), .valid_in_4(valid_in_164), .pxl_in_4(pxl_in_164), .valid_in_5(valid_in_165), .pxl_in_5(pxl_in_165), .valid_in_6(valid_in_166), .pxl_in_6(pxl_in_166), .valid_in_7(valid_in_167), .pxl_in_7(pxl_in_167), .valid_in_8(valid_in_168), .pxl_in_8(pxl_in_168), .valid_in_9(valid_in_169), .pxl_in_9(pxl_in_169), .valid_in_10(valid_in_170), .pxl_in_10(pxl_in_170), .valid_in_11(valid_in_171), .pxl_in_11(pxl_in_171), .valid_in_12(valid_in_172), .pxl_in_12(pxl_in_172), .valid_in_13(valid_in_173), .pxl_in_13(pxl_in_173), .valid_in_14(valid_in_174), .pxl_in_14(pxl_in_174), .valid_in_15(valid_in_175), .pxl_in_15(pxl_in_175), .valid_in_16(valid_in_176), .pxl_in_16(pxl_in_176), .valid_in_17(valid_in_177), .pxl_in_17(pxl_in_177), .valid_in_18(valid_in_178), .pxl_in_18(pxl_in_178), .valid_in_19(valid_in_179), .pxl_in_19(pxl_in_179), .valid_in_20(valid_in_180), .pxl_in_20(pxl_in_180), .valid_in_21(valid_in_181), .pxl_in_21(pxl_in_181), .valid_in_22(valid_in_182), .pxl_in_22(pxl_in_182), .valid_in_23(valid_in_183), .pxl_in_23(pxl_in_183), .valid_in_24(valid_in_184), .pxl_in_24(pxl_in_184), .valid_in_25(valid_in_185), .pxl_in_25(pxl_in_185), .valid_in_26(valid_in_186), .pxl_in_26(pxl_in_186), .valid_in_27(valid_in_187), .pxl_in_27(pxl_in_187), .valid_in_28(valid_in_188), .pxl_in_28(pxl_in_188), .valid_in_29(valid_in_189), .pxl_in_29(pxl_in_189), .valid_in_30(valid_in_190), .pxl_in_30(pxl_in_190), .valid_in_31(valid_in_191), .pxl_in_31(pxl_in_191), .valid_in_32(valid_in_192), .pxl_in_32(pxl_in_192), .pxl_out(pxl_out_6), .valid_out(valid_out_6) );

add_32layers#(D, DATA_WIDTH) x7(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_193), .pxl_in_1(pxl_in_193), .valid_in_2(valid_in_194), .pxl_in_2(pxl_in_194), .valid_in_3(valid_in_195), .pxl_in_3(pxl_in_195), .valid_in_4(valid_in_196), .pxl_in_4(pxl_in_196), .valid_in_5(valid_in_197), .pxl_in_5(pxl_in_197), .valid_in_6(valid_in_198), .pxl_in_6(pxl_in_198), .valid_in_7(valid_in_199), .pxl_in_7(pxl_in_199), .valid_in_8(valid_in_200), .pxl_in_8(pxl_in_200), .valid_in_9(valid_in_201), .pxl_in_9(pxl_in_201), .valid_in_10(valid_in_202), .pxl_in_10(pxl_in_202), .valid_in_11(valid_in_203), .pxl_in_11(pxl_in_203), .valid_in_12(valid_in_204), .pxl_in_12(pxl_in_204), .valid_in_13(valid_in_205), .pxl_in_13(pxl_in_205), .valid_in_14(valid_in_206), .pxl_in_14(pxl_in_206), .valid_in_15(valid_in_207), .pxl_in_15(pxl_in_207), .valid_in_16(valid_in_208), .pxl_in_16(pxl_in_208), .valid_in_17(valid_in_209), .pxl_in_17(pxl_in_209), .valid_in_18(valid_in_210), .pxl_in_18(pxl_in_210), .valid_in_19(valid_in_211), .pxl_in_19(pxl_in_211), .valid_in_20(valid_in_212), .pxl_in_20(pxl_in_212), .valid_in_21(valid_in_213), .pxl_in_21(pxl_in_213), .valid_in_22(valid_in_214), .pxl_in_22(pxl_in_214), .valid_in_23(valid_in_215), .pxl_in_23(pxl_in_215), .valid_in_24(valid_in_216), .pxl_in_24(pxl_in_216), .valid_in_25(valid_in_217), .pxl_in_25(pxl_in_217), .valid_in_26(valid_in_218), .pxl_in_26(pxl_in_218), .valid_in_27(valid_in_219), .pxl_in_27(pxl_in_219), .valid_in_28(valid_in_220), .pxl_in_28(pxl_in_220), .valid_in_29(valid_in_221), .pxl_in_29(pxl_in_221), .valid_in_30(valid_in_222), .pxl_in_30(pxl_in_222), .valid_in_31(valid_in_223), .pxl_in_31(pxl_in_223), .valid_in_32(valid_in_224), .pxl_in_32(pxl_in_224), .pxl_out(pxl_out_7), .valid_out(valid_out_7) );

add_32layers#(D, DATA_WIDTH) x8(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_225), .pxl_in_1(pxl_in_225), .valid_in_2(valid_in_226), .pxl_in_2(pxl_in_226), .valid_in_3(valid_in_227), .pxl_in_3(pxl_in_227), .valid_in_4(valid_in_228), .pxl_in_4(pxl_in_228), .valid_in_5(valid_in_229), .pxl_in_5(pxl_in_229), .valid_in_6(valid_in_230), .pxl_in_6(pxl_in_230), .valid_in_7(valid_in_231), .pxl_in_7(pxl_in_231), .valid_in_8(valid_in_232), .pxl_in_8(pxl_in_232), .valid_in_9(valid_in_233), .pxl_in_9(pxl_in_233), .valid_in_10(valid_in_234), .pxl_in_10(pxl_in_234), .valid_in_11(valid_in_235), .pxl_in_11(pxl_in_235), .valid_in_12(valid_in_236), .pxl_in_12(pxl_in_236), .valid_in_13(valid_in_237), .pxl_in_13(pxl_in_237), .valid_in_14(valid_in_238), .pxl_in_14(pxl_in_238), .valid_in_15(valid_in_239), .pxl_in_15(pxl_in_239), .valid_in_16(valid_in_240), .pxl_in_16(pxl_in_240), .valid_in_17(valid_in_241), .pxl_in_17(pxl_in_241), .valid_in_18(valid_in_242), .pxl_in_18(pxl_in_242), .valid_in_19(valid_in_243), .pxl_in_19(pxl_in_243), .valid_in_20(valid_in_244), .pxl_in_20(pxl_in_244), .valid_in_21(valid_in_245), .pxl_in_21(pxl_in_245), .valid_in_22(valid_in_246), .pxl_in_22(pxl_in_246), .valid_in_23(valid_in_247), .pxl_in_23(pxl_in_247), .valid_in_24(valid_in_248), .pxl_in_24(pxl_in_248), .valid_in_25(valid_in_249), .pxl_in_25(pxl_in_249), .valid_in_26(valid_in_250), .pxl_in_26(pxl_in_250), .valid_in_27(valid_in_251), .pxl_in_27(pxl_in_251), .valid_in_28(valid_in_252), .pxl_in_28(pxl_in_252), .valid_in_29(valid_in_253), .pxl_in_29(pxl_in_253), .valid_in_30(valid_in_254), .pxl_in_30(pxl_in_254), .valid_in_31(valid_in_255), .pxl_in_31(pxl_in_255), .valid_in_32(valid_in_256), .pxl_in_32(pxl_in_256), .pxl_out(pxl_out_8), .valid_out(valid_out_8) );

add_32layers#(D, DATA_WIDTH) x9(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_257), .pxl_in_1(pxl_in_257), .valid_in_2(valid_in_258), .pxl_in_2(pxl_in_258), .valid_in_3(valid_in_259), .pxl_in_3(pxl_in_259), .valid_in_4(valid_in_260), .pxl_in_4(pxl_in_260), .valid_in_5(valid_in_261), .pxl_in_5(pxl_in_261), .valid_in_6(valid_in_262), .pxl_in_6(pxl_in_262), .valid_in_7(valid_in_263), .pxl_in_7(pxl_in_263), .valid_in_8(valid_in_264), .pxl_in_8(pxl_in_264), .valid_in_9(valid_in_265), .pxl_in_9(pxl_in_265), .valid_in_10(valid_in_266), .pxl_in_10(pxl_in_266), .valid_in_11(valid_in_267), .pxl_in_11(pxl_in_267), .valid_in_12(valid_in_268), .pxl_in_12(pxl_in_268), .valid_in_13(valid_in_269), .pxl_in_13(pxl_in_269), .valid_in_14(valid_in_270), .pxl_in_14(pxl_in_270), .valid_in_15(valid_in_271), .pxl_in_15(pxl_in_271), .valid_in_16(valid_in_272), .pxl_in_16(pxl_in_272), .valid_in_17(valid_in_273), .pxl_in_17(pxl_in_273), .valid_in_18(valid_in_274), .pxl_in_18(pxl_in_274), .valid_in_19(valid_in_275), .pxl_in_19(pxl_in_275), .valid_in_20(valid_in_276), .pxl_in_20(pxl_in_276), .valid_in_21(valid_in_277), .pxl_in_21(pxl_in_277), .valid_in_22(valid_in_278), .pxl_in_22(pxl_in_278), .valid_in_23(valid_in_279), .pxl_in_23(pxl_in_279), .valid_in_24(valid_in_280), .pxl_in_24(pxl_in_280), .valid_in_25(valid_in_281), .pxl_in_25(pxl_in_281), .valid_in_26(valid_in_282), .pxl_in_26(pxl_in_282), .valid_in_27(valid_in_283), .pxl_in_27(pxl_in_283), .valid_in_28(valid_in_284), .pxl_in_28(pxl_in_284), .valid_in_29(valid_in_285), .pxl_in_29(pxl_in_285), .valid_in_30(valid_in_286), .pxl_in_30(pxl_in_286), .valid_in_31(valid_in_287), .pxl_in_31(pxl_in_287), .valid_in_32(valid_in_288), .pxl_in_32(pxl_in_288), .pxl_out(pxl_out_9), .valid_out(valid_out_9) );

add_32layers#(D, DATA_WIDTH) x10(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_289), .pxl_in_1(pxl_in_289), .valid_in_2(valid_in_290), .pxl_in_2(pxl_in_290), .valid_in_3(valid_in_291), .pxl_in_3(pxl_in_291), .valid_in_4(valid_in_292), .pxl_in_4(pxl_in_292), .valid_in_5(valid_in_293), .pxl_in_5(pxl_in_293), .valid_in_6(valid_in_294), .pxl_in_6(pxl_in_294), .valid_in_7(valid_in_295), .pxl_in_7(pxl_in_295), .valid_in_8(valid_in_296), .pxl_in_8(pxl_in_296), .valid_in_9(valid_in_297), .pxl_in_9(pxl_in_297), .valid_in_10(valid_in_298), .pxl_in_10(pxl_in_298), .valid_in_11(valid_in_299), .pxl_in_11(pxl_in_299), .valid_in_12(valid_in_300), .pxl_in_12(pxl_in_300), .valid_in_13(valid_in_301), .pxl_in_13(pxl_in_301), .valid_in_14(valid_in_302), .pxl_in_14(pxl_in_302), .valid_in_15(valid_in_303), .pxl_in_15(pxl_in_303), .valid_in_16(valid_in_304), .pxl_in_16(pxl_in_304), .valid_in_17(valid_in_305), .pxl_in_17(pxl_in_305), .valid_in_18(valid_in_306), .pxl_in_18(pxl_in_306), .valid_in_19(valid_in_307), .pxl_in_19(pxl_in_307), .valid_in_20(valid_in_308), .pxl_in_20(pxl_in_308), .valid_in_21(valid_in_309), .pxl_in_21(pxl_in_309), .valid_in_22(valid_in_310), .pxl_in_22(pxl_in_310), .valid_in_23(valid_in_311), .pxl_in_23(pxl_in_311), .valid_in_24(valid_in_312), .pxl_in_24(pxl_in_312), .valid_in_25(valid_in_313), .pxl_in_25(pxl_in_313), .valid_in_26(valid_in_314), .pxl_in_26(pxl_in_314), .valid_in_27(valid_in_315), .pxl_in_27(pxl_in_315), .valid_in_28(valid_in_316), .pxl_in_28(pxl_in_316), .valid_in_29(valid_in_317), .pxl_in_29(pxl_in_317), .valid_in_30(valid_in_318), .pxl_in_30(pxl_in_318), .valid_in_31(valid_in_319), .pxl_in_31(pxl_in_319), .valid_in_32(valid_in_320), .pxl_in_32(pxl_in_320), .pxl_out(pxl_out_10), .valid_out(valid_out_10) );

add_32layers#(D, DATA_WIDTH) x11(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_321), .pxl_in_1(pxl_in_321), .valid_in_2(valid_in_322), .pxl_in_2(pxl_in_322), .valid_in_3(valid_in_323), .pxl_in_3(pxl_in_323), .valid_in_4(valid_in_324), .pxl_in_4(pxl_in_324), .valid_in_5(valid_in_325), .pxl_in_5(pxl_in_325), .valid_in_6(valid_in_326), .pxl_in_6(pxl_in_326), .valid_in_7(valid_in_327), .pxl_in_7(pxl_in_327), .valid_in_8(valid_in_328), .pxl_in_8(pxl_in_328), .valid_in_9(valid_in_329), .pxl_in_9(pxl_in_329), .valid_in_10(valid_in_330), .pxl_in_10(pxl_in_330), .valid_in_11(valid_in_331), .pxl_in_11(pxl_in_331), .valid_in_12(valid_in_332), .pxl_in_12(pxl_in_332), .valid_in_13(valid_in_333), .pxl_in_13(pxl_in_333), .valid_in_14(valid_in_334), .pxl_in_14(pxl_in_334), .valid_in_15(valid_in_335), .pxl_in_15(pxl_in_335), .valid_in_16(valid_in_336), .pxl_in_16(pxl_in_336), .valid_in_17(valid_in_337), .pxl_in_17(pxl_in_337), .valid_in_18(valid_in_338), .pxl_in_18(pxl_in_338), .valid_in_19(valid_in_339), .pxl_in_19(pxl_in_339), .valid_in_20(valid_in_340), .pxl_in_20(pxl_in_340), .valid_in_21(valid_in_341), .pxl_in_21(pxl_in_341), .valid_in_22(valid_in_342), .pxl_in_22(pxl_in_342), .valid_in_23(valid_in_343), .pxl_in_23(pxl_in_343), .valid_in_24(valid_in_344), .pxl_in_24(pxl_in_344), .valid_in_25(valid_in_345), .pxl_in_25(pxl_in_345), .valid_in_26(valid_in_346), .pxl_in_26(pxl_in_346), .valid_in_27(valid_in_347), .pxl_in_27(pxl_in_347), .valid_in_28(valid_in_348), .pxl_in_28(pxl_in_348), .valid_in_29(valid_in_349), .pxl_in_29(pxl_in_349), .valid_in_30(valid_in_350), .pxl_in_30(pxl_in_350), .valid_in_31(valid_in_351), .pxl_in_31(pxl_in_351), .valid_in_32(valid_in_352), .pxl_in_32(pxl_in_352), .pxl_out(pxl_out_11), .valid_out(valid_out_11) );

add_32layers#(D, DATA_WIDTH) x12(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_353), .pxl_in_1(pxl_in_353), .valid_in_2(valid_in_354), .pxl_in_2(pxl_in_354), .valid_in_3(valid_in_355), .pxl_in_3(pxl_in_355), .valid_in_4(valid_in_356), .pxl_in_4(pxl_in_356), .valid_in_5(valid_in_357), .pxl_in_5(pxl_in_357), .valid_in_6(valid_in_358), .pxl_in_6(pxl_in_358), .valid_in_7(valid_in_359), .pxl_in_7(pxl_in_359), .valid_in_8(valid_in_360), .pxl_in_8(pxl_in_360), .valid_in_9(valid_in_361), .pxl_in_9(pxl_in_361), .valid_in_10(valid_in_362), .pxl_in_10(pxl_in_362), .valid_in_11(valid_in_363), .pxl_in_11(pxl_in_363), .valid_in_12(valid_in_364), .pxl_in_12(pxl_in_364), .valid_in_13(valid_in_365), .pxl_in_13(pxl_in_365), .valid_in_14(valid_in_366), .pxl_in_14(pxl_in_366), .valid_in_15(valid_in_367), .pxl_in_15(pxl_in_367), .valid_in_16(valid_in_368), .pxl_in_16(pxl_in_368), .valid_in_17(valid_in_369), .pxl_in_17(pxl_in_369), .valid_in_18(valid_in_370), .pxl_in_18(pxl_in_370), .valid_in_19(valid_in_371), .pxl_in_19(pxl_in_371), .valid_in_20(valid_in_372), .pxl_in_20(pxl_in_372), .valid_in_21(valid_in_373), .pxl_in_21(pxl_in_373), .valid_in_22(valid_in_374), .pxl_in_22(pxl_in_374), .valid_in_23(valid_in_375), .pxl_in_23(pxl_in_375), .valid_in_24(valid_in_376), .pxl_in_24(pxl_in_376), .valid_in_25(valid_in_377), .pxl_in_25(pxl_in_377), .valid_in_26(valid_in_378), .pxl_in_26(pxl_in_378), .valid_in_27(valid_in_379), .pxl_in_27(pxl_in_379), .valid_in_28(valid_in_380), .pxl_in_28(pxl_in_380), .valid_in_29(valid_in_381), .pxl_in_29(pxl_in_381), .valid_in_30(valid_in_382), .pxl_in_30(pxl_in_382), .valid_in_31(valid_in_383), .pxl_in_31(pxl_in_383), .valid_in_32(valid_in_384), .pxl_in_32(pxl_in_384), .pxl_out(pxl_out_12), .valid_out(valid_out_12) );

add_32layers#(D, DATA_WIDTH) x13(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_385), .pxl_in_1(pxl_in_385), .valid_in_2(valid_in_386), .pxl_in_2(pxl_in_386), .valid_in_3(valid_in_387), .pxl_in_3(pxl_in_387), .valid_in_4(valid_in_388), .pxl_in_4(pxl_in_388), .valid_in_5(valid_in_389), .pxl_in_5(pxl_in_389), .valid_in_6(valid_in_390), .pxl_in_6(pxl_in_390), .valid_in_7(valid_in_391), .pxl_in_7(pxl_in_391), .valid_in_8(valid_in_392), .pxl_in_8(pxl_in_392), .valid_in_9(valid_in_393), .pxl_in_9(pxl_in_393), .valid_in_10(valid_in_394), .pxl_in_10(pxl_in_394), .valid_in_11(valid_in_395), .pxl_in_11(pxl_in_395), .valid_in_12(valid_in_396), .pxl_in_12(pxl_in_396), .valid_in_13(valid_in_397), .pxl_in_13(pxl_in_397), .valid_in_14(valid_in_398), .pxl_in_14(pxl_in_398), .valid_in_15(valid_in_399), .pxl_in_15(pxl_in_399), .valid_in_16(valid_in_400), .pxl_in_16(pxl_in_400), .valid_in_17(valid_in_401), .pxl_in_17(pxl_in_401), .valid_in_18(valid_in_402), .pxl_in_18(pxl_in_402), .valid_in_19(valid_in_403), .pxl_in_19(pxl_in_403), .valid_in_20(valid_in_404), .pxl_in_20(pxl_in_404), .valid_in_21(valid_in_405), .pxl_in_21(pxl_in_405), .valid_in_22(valid_in_406), .pxl_in_22(pxl_in_406), .valid_in_23(valid_in_407), .pxl_in_23(pxl_in_407), .valid_in_24(valid_in_408), .pxl_in_24(pxl_in_408), .valid_in_25(valid_in_409), .pxl_in_25(pxl_in_409), .valid_in_26(valid_in_410), .pxl_in_26(pxl_in_410), .valid_in_27(valid_in_411), .pxl_in_27(pxl_in_411), .valid_in_28(valid_in_412), .pxl_in_28(pxl_in_412), .valid_in_29(valid_in_413), .pxl_in_29(pxl_in_413), .valid_in_30(valid_in_414), .pxl_in_30(pxl_in_414), .valid_in_31(valid_in_415), .pxl_in_31(pxl_in_415), .valid_in_32(valid_in_416), .pxl_in_32(pxl_in_416), .pxl_out(pxl_out_13), .valid_out(valid_out_13) );

add_32layers#(D, DATA_WIDTH) x14(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_417), .pxl_in_1(pxl_in_417), .valid_in_2(valid_in_418), .pxl_in_2(pxl_in_418), .valid_in_3(valid_in_419), .pxl_in_3(pxl_in_419), .valid_in_4(valid_in_420), .pxl_in_4(pxl_in_420), .valid_in_5(valid_in_421), .pxl_in_5(pxl_in_421), .valid_in_6(valid_in_422), .pxl_in_6(pxl_in_422), .valid_in_7(valid_in_423), .pxl_in_7(pxl_in_423), .valid_in_8(valid_in_424), .pxl_in_8(pxl_in_424), .valid_in_9(valid_in_425), .pxl_in_9(pxl_in_425), .valid_in_10(valid_in_426), .pxl_in_10(pxl_in_426), .valid_in_11(valid_in_427), .pxl_in_11(pxl_in_427), .valid_in_12(valid_in_428), .pxl_in_12(pxl_in_428), .valid_in_13(valid_in_429), .pxl_in_13(pxl_in_429), .valid_in_14(valid_in_430), .pxl_in_14(pxl_in_430), .valid_in_15(valid_in_431), .pxl_in_15(pxl_in_431), .valid_in_16(valid_in_432), .pxl_in_16(pxl_in_432), .valid_in_17(valid_in_433), .pxl_in_17(pxl_in_433), .valid_in_18(valid_in_434), .pxl_in_18(pxl_in_434), .valid_in_19(valid_in_435), .pxl_in_19(pxl_in_435), .valid_in_20(valid_in_436), .pxl_in_20(pxl_in_436), .valid_in_21(valid_in_437), .pxl_in_21(pxl_in_437), .valid_in_22(valid_in_438), .pxl_in_22(pxl_in_438), .valid_in_23(valid_in_439), .pxl_in_23(pxl_in_439), .valid_in_24(valid_in_440), .pxl_in_24(pxl_in_440), .valid_in_25(valid_in_441), .pxl_in_25(pxl_in_441), .valid_in_26(valid_in_442), .pxl_in_26(pxl_in_442), .valid_in_27(valid_in_443), .pxl_in_27(pxl_in_443), .valid_in_28(valid_in_444), .pxl_in_28(pxl_in_444), .valid_in_29(valid_in_445), .pxl_in_29(pxl_in_445), .valid_in_30(valid_in_446), .pxl_in_30(pxl_in_446), .valid_in_31(valid_in_447), .pxl_in_31(pxl_in_447), .valid_in_32(valid_in_448), .pxl_in_32(pxl_in_448), .pxl_out(pxl_out_14), .valid_out(valid_out_14) );

add_32layers#(D, DATA_WIDTH) x15(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_449), .pxl_in_1(pxl_in_449), .valid_in_2(valid_in_450), .pxl_in_2(pxl_in_450), .valid_in_3(valid_in_451), .pxl_in_3(pxl_in_451), .valid_in_4(valid_in_452), .pxl_in_4(pxl_in_452), .valid_in_5(valid_in_453), .pxl_in_5(pxl_in_453), .valid_in_6(valid_in_454), .pxl_in_6(pxl_in_454), .valid_in_7(valid_in_455), .pxl_in_7(pxl_in_455), .valid_in_8(valid_in_456), .pxl_in_8(pxl_in_456), .valid_in_9(valid_in_457), .pxl_in_9(pxl_in_457), .valid_in_10(valid_in_458), .pxl_in_10(pxl_in_458), .valid_in_11(valid_in_459), .pxl_in_11(pxl_in_459), .valid_in_12(valid_in_460), .pxl_in_12(pxl_in_460), .valid_in_13(valid_in_461), .pxl_in_13(pxl_in_461), .valid_in_14(valid_in_462), .pxl_in_14(pxl_in_462), .valid_in_15(valid_in_463), .pxl_in_15(pxl_in_463), .valid_in_16(valid_in_464), .pxl_in_16(pxl_in_464), .valid_in_17(valid_in_465), .pxl_in_17(pxl_in_465), .valid_in_18(valid_in_466), .pxl_in_18(pxl_in_466), .valid_in_19(valid_in_467), .pxl_in_19(pxl_in_467), .valid_in_20(valid_in_468), .pxl_in_20(pxl_in_468), .valid_in_21(valid_in_469), .pxl_in_21(pxl_in_469), .valid_in_22(valid_in_470), .pxl_in_22(pxl_in_470), .valid_in_23(valid_in_471), .pxl_in_23(pxl_in_471), .valid_in_24(valid_in_472), .pxl_in_24(pxl_in_472), .valid_in_25(valid_in_473), .pxl_in_25(pxl_in_473), .valid_in_26(valid_in_474), .pxl_in_26(pxl_in_474), .valid_in_27(valid_in_475), .pxl_in_27(pxl_in_475), .valid_in_28(valid_in_476), .pxl_in_28(pxl_in_476), .valid_in_29(valid_in_477), .pxl_in_29(pxl_in_477), .valid_in_30(valid_in_478), .pxl_in_30(pxl_in_478), .valid_in_31(valid_in_479), .pxl_in_31(pxl_in_479), .valid_in_32(valid_in_480), .pxl_in_32(pxl_in_480), .pxl_out(pxl_out_15), .valid_out(valid_out_15) );

add_32layers#(D, DATA_WIDTH) x16(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_481), .pxl_in_1(pxl_in_481), .valid_in_2(valid_in_482), .pxl_in_2(pxl_in_482), .valid_in_3(valid_in_483), .pxl_in_3(pxl_in_483), .valid_in_4(valid_in_484), .pxl_in_4(pxl_in_484), .valid_in_5(valid_in_485), .pxl_in_5(pxl_in_485), .valid_in_6(valid_in_486), .pxl_in_6(pxl_in_486), .valid_in_7(valid_in_487), .pxl_in_7(pxl_in_487), .valid_in_8(valid_in_488), .pxl_in_8(pxl_in_488), .valid_in_9(valid_in_489), .pxl_in_9(pxl_in_489), .valid_in_10(valid_in_490), .pxl_in_10(pxl_in_490), .valid_in_11(valid_in_491), .pxl_in_11(pxl_in_491), .valid_in_12(valid_in_492), .pxl_in_12(pxl_in_492), .valid_in_13(valid_in_493), .pxl_in_13(pxl_in_493), .valid_in_14(valid_in_494), .pxl_in_14(pxl_in_494), .valid_in_15(valid_in_495), .pxl_in_15(pxl_in_495), .valid_in_16(valid_in_496), .pxl_in_16(pxl_in_496), .valid_in_17(valid_in_497), .pxl_in_17(pxl_in_497), .valid_in_18(valid_in_498), .pxl_in_18(pxl_in_498), .valid_in_19(valid_in_499), .pxl_in_19(pxl_in_499), .valid_in_20(valid_in_500), .pxl_in_20(pxl_in_500), .valid_in_21(valid_in_501), .pxl_in_21(pxl_in_501), .valid_in_22(valid_in_502), .pxl_in_22(pxl_in_502), .valid_in_23(valid_in_503), .pxl_in_23(pxl_in_503), .valid_in_24(valid_in_504), .pxl_in_24(pxl_in_504), .valid_in_25(valid_in_505), .pxl_in_25(pxl_in_505), .valid_in_26(valid_in_506), .pxl_in_26(pxl_in_506), .valid_in_27(valid_in_507), .pxl_in_27(pxl_in_507), .valid_in_28(valid_in_508), .pxl_in_28(pxl_in_508), .valid_in_29(valid_in_509), .pxl_in_29(pxl_in_509), .valid_in_30(valid_in_510), .pxl_in_30(pxl_in_510), .valid_in_31(valid_in_511), .pxl_in_31(pxl_in_511), .valid_in_32(valid_in_512), .pxl_in_32(pxl_in_512), .pxl_out(pxl_out_16), .valid_out(valid_out_16) );

add_32layers#(D, DATA_WIDTH) x17(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_513), .pxl_in_1(pxl_in_513), .valid_in_2(valid_in_514), .pxl_in_2(pxl_in_514), .valid_in_3(valid_in_515), .pxl_in_3(pxl_in_515), .valid_in_4(valid_in_516), .pxl_in_4(pxl_in_516), .valid_in_5(valid_in_517), .pxl_in_5(pxl_in_517), .valid_in_6(valid_in_518), .pxl_in_6(pxl_in_518), .valid_in_7(valid_in_519), .pxl_in_7(pxl_in_519), .valid_in_8(valid_in_520), .pxl_in_8(pxl_in_520), .valid_in_9(valid_in_521), .pxl_in_9(pxl_in_521), .valid_in_10(valid_in_522), .pxl_in_10(pxl_in_522), .valid_in_11(valid_in_523), .pxl_in_11(pxl_in_523), .valid_in_12(valid_in_524), .pxl_in_12(pxl_in_524), .valid_in_13(valid_in_525), .pxl_in_13(pxl_in_525), .valid_in_14(valid_in_526), .pxl_in_14(pxl_in_526), .valid_in_15(valid_in_527), .pxl_in_15(pxl_in_527), .valid_in_16(valid_in_528), .pxl_in_16(pxl_in_528), .valid_in_17(valid_in_529), .pxl_in_17(pxl_in_529), .valid_in_18(valid_in_530), .pxl_in_18(pxl_in_530), .valid_in_19(valid_in_531), .pxl_in_19(pxl_in_531), .valid_in_20(valid_in_532), .pxl_in_20(pxl_in_532), .valid_in_21(valid_in_533), .pxl_in_21(pxl_in_533), .valid_in_22(valid_in_534), .pxl_in_22(pxl_in_534), .valid_in_23(valid_in_535), .pxl_in_23(pxl_in_535), .valid_in_24(valid_in_536), .pxl_in_24(pxl_in_536), .valid_in_25(valid_in_537), .pxl_in_25(pxl_in_537), .valid_in_26(valid_in_538), .pxl_in_26(pxl_in_538), .valid_in_27(valid_in_539), .pxl_in_27(pxl_in_539), .valid_in_28(valid_in_540), .pxl_in_28(pxl_in_540), .valid_in_29(valid_in_541), .pxl_in_29(pxl_in_541), .valid_in_30(valid_in_542), .pxl_in_30(pxl_in_542), .valid_in_31(valid_in_543), .pxl_in_31(pxl_in_543), .valid_in_32(valid_in_544), .pxl_in_32(pxl_in_544), .pxl_out(pxl_out_17), .valid_out(valid_out_17) );

add_32layers#(D, DATA_WIDTH) x18(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_545), .pxl_in_1(pxl_in_545), .valid_in_2(valid_in_546), .pxl_in_2(pxl_in_546), .valid_in_3(valid_in_547), .pxl_in_3(pxl_in_547), .valid_in_4(valid_in_548), .pxl_in_4(pxl_in_548), .valid_in_5(valid_in_549), .pxl_in_5(pxl_in_549), .valid_in_6(valid_in_550), .pxl_in_6(pxl_in_550), .valid_in_7(valid_in_551), .pxl_in_7(pxl_in_551), .valid_in_8(valid_in_552), .pxl_in_8(pxl_in_552), .valid_in_9(valid_in_553), .pxl_in_9(pxl_in_553), .valid_in_10(valid_in_554), .pxl_in_10(pxl_in_554), .valid_in_11(valid_in_555), .pxl_in_11(pxl_in_555), .valid_in_12(valid_in_556), .pxl_in_12(pxl_in_556), .valid_in_13(valid_in_557), .pxl_in_13(pxl_in_557), .valid_in_14(valid_in_558), .pxl_in_14(pxl_in_558), .valid_in_15(valid_in_559), .pxl_in_15(pxl_in_559), .valid_in_16(valid_in_560), .pxl_in_16(pxl_in_560), .valid_in_17(valid_in_561), .pxl_in_17(pxl_in_561), .valid_in_18(valid_in_562), .pxl_in_18(pxl_in_562), .valid_in_19(valid_in_563), .pxl_in_19(pxl_in_563), .valid_in_20(valid_in_564), .pxl_in_20(pxl_in_564), .valid_in_21(valid_in_565), .pxl_in_21(pxl_in_565), .valid_in_22(valid_in_566), .pxl_in_22(pxl_in_566), .valid_in_23(valid_in_567), .pxl_in_23(pxl_in_567), .valid_in_24(valid_in_568), .pxl_in_24(pxl_in_568), .valid_in_25(valid_in_569), .pxl_in_25(pxl_in_569), .valid_in_26(valid_in_570), .pxl_in_26(pxl_in_570), .valid_in_27(valid_in_571), .pxl_in_27(pxl_in_571), .valid_in_28(valid_in_572), .pxl_in_28(pxl_in_572), .valid_in_29(valid_in_573), .pxl_in_29(pxl_in_573), .valid_in_30(valid_in_574), .pxl_in_30(pxl_in_574), .valid_in_31(valid_in_575), .pxl_in_31(pxl_in_575), .valid_in_32(valid_in_576), .pxl_in_32(pxl_in_576), .pxl_out(pxl_out_18), .valid_out(valid_out_18) );

add_32layers#(D, DATA_WIDTH) x19(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_577), .pxl_in_1(pxl_in_577), .valid_in_2(valid_in_578), .pxl_in_2(pxl_in_578), .valid_in_3(valid_in_579), .pxl_in_3(pxl_in_579), .valid_in_4(valid_in_580), .pxl_in_4(pxl_in_580), .valid_in_5(valid_in_581), .pxl_in_5(pxl_in_581), .valid_in_6(valid_in_582), .pxl_in_6(pxl_in_582), .valid_in_7(valid_in_583), .pxl_in_7(pxl_in_583), .valid_in_8(valid_in_584), .pxl_in_8(pxl_in_584), .valid_in_9(valid_in_585), .pxl_in_9(pxl_in_585), .valid_in_10(valid_in_586), .pxl_in_10(pxl_in_586), .valid_in_11(valid_in_587), .pxl_in_11(pxl_in_587), .valid_in_12(valid_in_588), .pxl_in_12(pxl_in_588), .valid_in_13(valid_in_589), .pxl_in_13(pxl_in_589), .valid_in_14(valid_in_590), .pxl_in_14(pxl_in_590), .valid_in_15(valid_in_591), .pxl_in_15(pxl_in_591), .valid_in_16(valid_in_592), .pxl_in_16(pxl_in_592), .valid_in_17(valid_in_593), .pxl_in_17(pxl_in_593), .valid_in_18(valid_in_594), .pxl_in_18(pxl_in_594), .valid_in_19(valid_in_595), .pxl_in_19(pxl_in_595), .valid_in_20(valid_in_596), .pxl_in_20(pxl_in_596), .valid_in_21(valid_in_597), .pxl_in_21(pxl_in_597), .valid_in_22(valid_in_598), .pxl_in_22(pxl_in_598), .valid_in_23(valid_in_599), .pxl_in_23(pxl_in_599), .valid_in_24(valid_in_600), .pxl_in_24(pxl_in_600), .valid_in_25(valid_in_601), .pxl_in_25(pxl_in_601), .valid_in_26(valid_in_602), .pxl_in_26(pxl_in_602), .valid_in_27(valid_in_603), .pxl_in_27(pxl_in_603), .valid_in_28(valid_in_604), .pxl_in_28(pxl_in_604), .valid_in_29(valid_in_605), .pxl_in_29(pxl_in_605), .valid_in_30(valid_in_606), .pxl_in_30(pxl_in_606), .valid_in_31(valid_in_607), .pxl_in_31(pxl_in_607), .valid_in_32(valid_in_608), .pxl_in_32(pxl_in_608), .pxl_out(pxl_out_19), .valid_out(valid_out_19) );

add_32layers#(D, DATA_WIDTH) x20(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_609), .pxl_in_1(pxl_in_609), .valid_in_2(valid_in_610), .pxl_in_2(pxl_in_610), .valid_in_3(valid_in_611), .pxl_in_3(pxl_in_611), .valid_in_4(valid_in_612), .pxl_in_4(pxl_in_612), .valid_in_5(valid_in_613), .pxl_in_5(pxl_in_613), .valid_in_6(valid_in_614), .pxl_in_6(pxl_in_614), .valid_in_7(valid_in_615), .pxl_in_7(pxl_in_615), .valid_in_8(valid_in_616), .pxl_in_8(pxl_in_616), .valid_in_9(valid_in_617), .pxl_in_9(pxl_in_617), .valid_in_10(valid_in_618), .pxl_in_10(pxl_in_618), .valid_in_11(valid_in_619), .pxl_in_11(pxl_in_619), .valid_in_12(valid_in_620), .pxl_in_12(pxl_in_620), .valid_in_13(valid_in_621), .pxl_in_13(pxl_in_621), .valid_in_14(valid_in_622), .pxl_in_14(pxl_in_622), .valid_in_15(valid_in_623), .pxl_in_15(pxl_in_623), .valid_in_16(valid_in_624), .pxl_in_16(pxl_in_624), .valid_in_17(valid_in_625), .pxl_in_17(pxl_in_625), .valid_in_18(valid_in_626), .pxl_in_18(pxl_in_626), .valid_in_19(valid_in_627), .pxl_in_19(pxl_in_627), .valid_in_20(valid_in_628), .pxl_in_20(pxl_in_628), .valid_in_21(valid_in_629), .pxl_in_21(pxl_in_629), .valid_in_22(valid_in_630), .pxl_in_22(pxl_in_630), .valid_in_23(valid_in_631), .pxl_in_23(pxl_in_631), .valid_in_24(valid_in_632), .pxl_in_24(pxl_in_632), .valid_in_25(valid_in_633), .pxl_in_25(pxl_in_633), .valid_in_26(valid_in_634), .pxl_in_26(pxl_in_634), .valid_in_27(valid_in_635), .pxl_in_27(pxl_in_635), .valid_in_28(valid_in_636), .pxl_in_28(pxl_in_636), .valid_in_29(valid_in_637), .pxl_in_29(pxl_in_637), .valid_in_30(valid_in_638), .pxl_in_30(pxl_in_638), .valid_in_31(valid_in_639), .pxl_in_31(pxl_in_639), .valid_in_32(valid_in_640), .pxl_in_32(pxl_in_640), .pxl_out(pxl_out_20), .valid_out(valid_out_20) );

add_32layers#(D, DATA_WIDTH) x21(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_641), .pxl_in_1(pxl_in_641), .valid_in_2(valid_in_642), .pxl_in_2(pxl_in_642), .valid_in_3(valid_in_643), .pxl_in_3(pxl_in_643), .valid_in_4(valid_in_644), .pxl_in_4(pxl_in_644), .valid_in_5(valid_in_645), .pxl_in_5(pxl_in_645), .valid_in_6(valid_in_646), .pxl_in_6(pxl_in_646), .valid_in_7(valid_in_647), .pxl_in_7(pxl_in_647), .valid_in_8(valid_in_648), .pxl_in_8(pxl_in_648), .valid_in_9(valid_in_649), .pxl_in_9(pxl_in_649), .valid_in_10(valid_in_650), .pxl_in_10(pxl_in_650), .valid_in_11(valid_in_651), .pxl_in_11(pxl_in_651), .valid_in_12(valid_in_652), .pxl_in_12(pxl_in_652), .valid_in_13(valid_in_653), .pxl_in_13(pxl_in_653), .valid_in_14(valid_in_654), .pxl_in_14(pxl_in_654), .valid_in_15(valid_in_655), .pxl_in_15(pxl_in_655), .valid_in_16(valid_in_656), .pxl_in_16(pxl_in_656), .valid_in_17(valid_in_657), .pxl_in_17(pxl_in_657), .valid_in_18(valid_in_658), .pxl_in_18(pxl_in_658), .valid_in_19(valid_in_659), .pxl_in_19(pxl_in_659), .valid_in_20(valid_in_660), .pxl_in_20(pxl_in_660), .valid_in_21(valid_in_661), .pxl_in_21(pxl_in_661), .valid_in_22(valid_in_662), .pxl_in_22(pxl_in_662), .valid_in_23(valid_in_663), .pxl_in_23(pxl_in_663), .valid_in_24(valid_in_664), .pxl_in_24(pxl_in_664), .valid_in_25(valid_in_665), .pxl_in_25(pxl_in_665), .valid_in_26(valid_in_666), .pxl_in_26(pxl_in_666), .valid_in_27(valid_in_667), .pxl_in_27(pxl_in_667), .valid_in_28(valid_in_668), .pxl_in_28(pxl_in_668), .valid_in_29(valid_in_669), .pxl_in_29(pxl_in_669), .valid_in_30(valid_in_670), .pxl_in_30(pxl_in_670), .valid_in_31(valid_in_671), .pxl_in_31(pxl_in_671), .valid_in_32(valid_in_672), .pxl_in_32(pxl_in_672), .pxl_out(pxl_out_21), .valid_out(valid_out_21) );

add_32layers#(D, DATA_WIDTH) x22(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_673), .pxl_in_1(pxl_in_673), .valid_in_2(valid_in_674), .pxl_in_2(pxl_in_674), .valid_in_3(valid_in_675), .pxl_in_3(pxl_in_675), .valid_in_4(valid_in_676), .pxl_in_4(pxl_in_676), .valid_in_5(valid_in_677), .pxl_in_5(pxl_in_677), .valid_in_6(valid_in_678), .pxl_in_6(pxl_in_678), .valid_in_7(valid_in_679), .pxl_in_7(pxl_in_679), .valid_in_8(valid_in_680), .pxl_in_8(pxl_in_680), .valid_in_9(valid_in_681), .pxl_in_9(pxl_in_681), .valid_in_10(valid_in_682), .pxl_in_10(pxl_in_682), .valid_in_11(valid_in_683), .pxl_in_11(pxl_in_683), .valid_in_12(valid_in_684), .pxl_in_12(pxl_in_684), .valid_in_13(valid_in_685), .pxl_in_13(pxl_in_685), .valid_in_14(valid_in_686), .pxl_in_14(pxl_in_686), .valid_in_15(valid_in_687), .pxl_in_15(pxl_in_687), .valid_in_16(valid_in_688), .pxl_in_16(pxl_in_688), .valid_in_17(valid_in_689), .pxl_in_17(pxl_in_689), .valid_in_18(valid_in_690), .pxl_in_18(pxl_in_690), .valid_in_19(valid_in_691), .pxl_in_19(pxl_in_691), .valid_in_20(valid_in_692), .pxl_in_20(pxl_in_692), .valid_in_21(valid_in_693), .pxl_in_21(pxl_in_693), .valid_in_22(valid_in_694), .pxl_in_22(pxl_in_694), .valid_in_23(valid_in_695), .pxl_in_23(pxl_in_695), .valid_in_24(valid_in_696), .pxl_in_24(pxl_in_696), .valid_in_25(valid_in_697), .pxl_in_25(pxl_in_697), .valid_in_26(valid_in_698), .pxl_in_26(pxl_in_698), .valid_in_27(valid_in_699), .pxl_in_27(pxl_in_699), .valid_in_28(valid_in_700), .pxl_in_28(pxl_in_700), .valid_in_29(valid_in_701), .pxl_in_29(pxl_in_701), .valid_in_30(valid_in_702), .pxl_in_30(pxl_in_702), .valid_in_31(valid_in_703), .pxl_in_31(pxl_in_703), .valid_in_32(valid_in_704), .pxl_in_32(pxl_in_704), .pxl_out(pxl_out_22), .valid_out(valid_out_22) );

add_32layers#(D, DATA_WIDTH) x23(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_705), .pxl_in_1(pxl_in_705), .valid_in_2(valid_in_706), .pxl_in_2(pxl_in_706), .valid_in_3(valid_in_707), .pxl_in_3(pxl_in_707), .valid_in_4(valid_in_708), .pxl_in_4(pxl_in_708), .valid_in_5(valid_in_709), .pxl_in_5(pxl_in_709), .valid_in_6(valid_in_710), .pxl_in_6(pxl_in_710), .valid_in_7(valid_in_711), .pxl_in_7(pxl_in_711), .valid_in_8(valid_in_712), .pxl_in_8(pxl_in_712), .valid_in_9(valid_in_713), .pxl_in_9(pxl_in_713), .valid_in_10(valid_in_714), .pxl_in_10(pxl_in_714), .valid_in_11(valid_in_715), .pxl_in_11(pxl_in_715), .valid_in_12(valid_in_716), .pxl_in_12(pxl_in_716), .valid_in_13(valid_in_717), .pxl_in_13(pxl_in_717), .valid_in_14(valid_in_718), .pxl_in_14(pxl_in_718), .valid_in_15(valid_in_719), .pxl_in_15(pxl_in_719), .valid_in_16(valid_in_720), .pxl_in_16(pxl_in_720), .valid_in_17(valid_in_721), .pxl_in_17(pxl_in_721), .valid_in_18(valid_in_722), .pxl_in_18(pxl_in_722), .valid_in_19(valid_in_723), .pxl_in_19(pxl_in_723), .valid_in_20(valid_in_724), .pxl_in_20(pxl_in_724), .valid_in_21(valid_in_725), .pxl_in_21(pxl_in_725), .valid_in_22(valid_in_726), .pxl_in_22(pxl_in_726), .valid_in_23(valid_in_727), .pxl_in_23(pxl_in_727), .valid_in_24(valid_in_728), .pxl_in_24(pxl_in_728), .valid_in_25(valid_in_729), .pxl_in_25(pxl_in_729), .valid_in_26(valid_in_730), .pxl_in_26(pxl_in_730), .valid_in_27(valid_in_731), .pxl_in_27(pxl_in_731), .valid_in_28(valid_in_732), .pxl_in_28(pxl_in_732), .valid_in_29(valid_in_733), .pxl_in_29(pxl_in_733), .valid_in_30(valid_in_734), .pxl_in_30(pxl_in_734), .valid_in_31(valid_in_735), .pxl_in_31(pxl_in_735), .valid_in_32(valid_in_736), .pxl_in_32(pxl_in_736), .pxl_out(pxl_out_23), .valid_out(valid_out_23) );

add_32layers#(D, DATA_WIDTH) x24(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_737), .pxl_in_1(pxl_in_737), .valid_in_2(valid_in_738), .pxl_in_2(pxl_in_738), .valid_in_3(valid_in_739), .pxl_in_3(pxl_in_739), .valid_in_4(valid_in_740), .pxl_in_4(pxl_in_740), .valid_in_5(valid_in_741), .pxl_in_5(pxl_in_741), .valid_in_6(valid_in_742), .pxl_in_6(pxl_in_742), .valid_in_7(valid_in_743), .pxl_in_7(pxl_in_743), .valid_in_8(valid_in_744), .pxl_in_8(pxl_in_744), .valid_in_9(valid_in_745), .pxl_in_9(pxl_in_745), .valid_in_10(valid_in_746), .pxl_in_10(pxl_in_746), .valid_in_11(valid_in_747), .pxl_in_11(pxl_in_747), .valid_in_12(valid_in_748), .pxl_in_12(pxl_in_748), .valid_in_13(valid_in_749), .pxl_in_13(pxl_in_749), .valid_in_14(valid_in_750), .pxl_in_14(pxl_in_750), .valid_in_15(valid_in_751), .pxl_in_15(pxl_in_751), .valid_in_16(valid_in_752), .pxl_in_16(pxl_in_752), .valid_in_17(valid_in_753), .pxl_in_17(pxl_in_753), .valid_in_18(valid_in_754), .pxl_in_18(pxl_in_754), .valid_in_19(valid_in_755), .pxl_in_19(pxl_in_755), .valid_in_20(valid_in_756), .pxl_in_20(pxl_in_756), .valid_in_21(valid_in_757), .pxl_in_21(pxl_in_757), .valid_in_22(valid_in_758), .pxl_in_22(pxl_in_758), .valid_in_23(valid_in_759), .pxl_in_23(pxl_in_759), .valid_in_24(valid_in_760), .pxl_in_24(pxl_in_760), .valid_in_25(valid_in_761), .pxl_in_25(pxl_in_761), .valid_in_26(valid_in_762), .pxl_in_26(pxl_in_762), .valid_in_27(valid_in_763), .pxl_in_27(pxl_in_763), .valid_in_28(valid_in_764), .pxl_in_28(pxl_in_764), .valid_in_29(valid_in_765), .pxl_in_29(pxl_in_765), .valid_in_30(valid_in_766), .pxl_in_30(pxl_in_766), .valid_in_31(valid_in_767), .pxl_in_31(pxl_in_767), .valid_in_32(valid_in_768), .pxl_in_32(pxl_in_768), .pxl_out(pxl_out_24), .valid_out(valid_out_24) );

add_32layers#(D, DATA_WIDTH) x25(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_769), .pxl_in_1(pxl_in_769), .valid_in_2(valid_in_770), .pxl_in_2(pxl_in_770), .valid_in_3(valid_in_771), .pxl_in_3(pxl_in_771), .valid_in_4(valid_in_772), .pxl_in_4(pxl_in_772), .valid_in_5(valid_in_773), .pxl_in_5(pxl_in_773), .valid_in_6(valid_in_774), .pxl_in_6(pxl_in_774), .valid_in_7(valid_in_775), .pxl_in_7(pxl_in_775), .valid_in_8(valid_in_776), .pxl_in_8(pxl_in_776), .valid_in_9(valid_in_777), .pxl_in_9(pxl_in_777), .valid_in_10(valid_in_778), .pxl_in_10(pxl_in_778), .valid_in_11(valid_in_779), .pxl_in_11(pxl_in_779), .valid_in_12(valid_in_780), .pxl_in_12(pxl_in_780), .valid_in_13(valid_in_781), .pxl_in_13(pxl_in_781), .valid_in_14(valid_in_782), .pxl_in_14(pxl_in_782), .valid_in_15(valid_in_783), .pxl_in_15(pxl_in_783), .valid_in_16(valid_in_784), .pxl_in_16(pxl_in_784), .valid_in_17(valid_in_785), .pxl_in_17(pxl_in_785), .valid_in_18(valid_in_786), .pxl_in_18(pxl_in_786), .valid_in_19(valid_in_787), .pxl_in_19(pxl_in_787), .valid_in_20(valid_in_788), .pxl_in_20(pxl_in_788), .valid_in_21(valid_in_789), .pxl_in_21(pxl_in_789), .valid_in_22(valid_in_790), .pxl_in_22(pxl_in_790), .valid_in_23(valid_in_791), .pxl_in_23(pxl_in_791), .valid_in_24(valid_in_792), .pxl_in_24(pxl_in_792), .valid_in_25(valid_in_793), .pxl_in_25(pxl_in_793), .valid_in_26(valid_in_794), .pxl_in_26(pxl_in_794), .valid_in_27(valid_in_795), .pxl_in_27(pxl_in_795), .valid_in_28(valid_in_796), .pxl_in_28(pxl_in_796), .valid_in_29(valid_in_797), .pxl_in_29(pxl_in_797), .valid_in_30(valid_in_798), .pxl_in_30(pxl_in_798), .valid_in_31(valid_in_799), .pxl_in_31(pxl_in_799), .valid_in_32(valid_in_800), .pxl_in_32(pxl_in_800), .pxl_out(pxl_out_25), .valid_out(valid_out_25) );

add_32layers#(D, DATA_WIDTH) x26(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_801), .pxl_in_1(pxl_in_801), .valid_in_2(valid_in_802), .pxl_in_2(pxl_in_802), .valid_in_3(valid_in_803), .pxl_in_3(pxl_in_803), .valid_in_4(valid_in_804), .pxl_in_4(pxl_in_804), .valid_in_5(valid_in_805), .pxl_in_5(pxl_in_805), .valid_in_6(valid_in_806), .pxl_in_6(pxl_in_806), .valid_in_7(valid_in_807), .pxl_in_7(pxl_in_807), .valid_in_8(valid_in_808), .pxl_in_8(pxl_in_808), .valid_in_9(valid_in_809), .pxl_in_9(pxl_in_809), .valid_in_10(valid_in_810), .pxl_in_10(pxl_in_810), .valid_in_11(valid_in_811), .pxl_in_11(pxl_in_811), .valid_in_12(valid_in_812), .pxl_in_12(pxl_in_812), .valid_in_13(valid_in_813), .pxl_in_13(pxl_in_813), .valid_in_14(valid_in_814), .pxl_in_14(pxl_in_814), .valid_in_15(valid_in_815), .pxl_in_15(pxl_in_815), .valid_in_16(valid_in_816), .pxl_in_16(pxl_in_816), .valid_in_17(valid_in_817), .pxl_in_17(pxl_in_817), .valid_in_18(valid_in_818), .pxl_in_18(pxl_in_818), .valid_in_19(valid_in_819), .pxl_in_19(pxl_in_819), .valid_in_20(valid_in_820), .pxl_in_20(pxl_in_820), .valid_in_21(valid_in_821), .pxl_in_21(pxl_in_821), .valid_in_22(valid_in_822), .pxl_in_22(pxl_in_822), .valid_in_23(valid_in_823), .pxl_in_23(pxl_in_823), .valid_in_24(valid_in_824), .pxl_in_24(pxl_in_824), .valid_in_25(valid_in_825), .pxl_in_25(pxl_in_825), .valid_in_26(valid_in_826), .pxl_in_26(pxl_in_826), .valid_in_27(valid_in_827), .pxl_in_27(pxl_in_827), .valid_in_28(valid_in_828), .pxl_in_28(pxl_in_828), .valid_in_29(valid_in_829), .pxl_in_29(pxl_in_829), .valid_in_30(valid_in_830), .pxl_in_30(pxl_in_830), .valid_in_31(valid_in_831), .pxl_in_31(pxl_in_831), .valid_in_32(valid_in_832), .pxl_in_32(pxl_in_832), .pxl_out(pxl_out_26), .valid_out(valid_out_26) );

add_32layers#(D, DATA_WIDTH) x27(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_833), .pxl_in_1(pxl_in_833), .valid_in_2(valid_in_834), .pxl_in_2(pxl_in_834), .valid_in_3(valid_in_835), .pxl_in_3(pxl_in_835), .valid_in_4(valid_in_836), .pxl_in_4(pxl_in_836), .valid_in_5(valid_in_837), .pxl_in_5(pxl_in_837), .valid_in_6(valid_in_838), .pxl_in_6(pxl_in_838), .valid_in_7(valid_in_839), .pxl_in_7(pxl_in_839), .valid_in_8(valid_in_840), .pxl_in_8(pxl_in_840), .valid_in_9(valid_in_841), .pxl_in_9(pxl_in_841), .valid_in_10(valid_in_842), .pxl_in_10(pxl_in_842), .valid_in_11(valid_in_843), .pxl_in_11(pxl_in_843), .valid_in_12(valid_in_844), .pxl_in_12(pxl_in_844), .valid_in_13(valid_in_845), .pxl_in_13(pxl_in_845), .valid_in_14(valid_in_846), .pxl_in_14(pxl_in_846), .valid_in_15(valid_in_847), .pxl_in_15(pxl_in_847), .valid_in_16(valid_in_848), .pxl_in_16(pxl_in_848), .valid_in_17(valid_in_849), .pxl_in_17(pxl_in_849), .valid_in_18(valid_in_850), .pxl_in_18(pxl_in_850), .valid_in_19(valid_in_851), .pxl_in_19(pxl_in_851), .valid_in_20(valid_in_852), .pxl_in_20(pxl_in_852), .valid_in_21(valid_in_853), .pxl_in_21(pxl_in_853), .valid_in_22(valid_in_854), .pxl_in_22(pxl_in_854), .valid_in_23(valid_in_855), .pxl_in_23(pxl_in_855), .valid_in_24(valid_in_856), .pxl_in_24(pxl_in_856), .valid_in_25(valid_in_857), .pxl_in_25(pxl_in_857), .valid_in_26(valid_in_858), .pxl_in_26(pxl_in_858), .valid_in_27(valid_in_859), .pxl_in_27(pxl_in_859), .valid_in_28(valid_in_860), .pxl_in_28(pxl_in_860), .valid_in_29(valid_in_861), .pxl_in_29(pxl_in_861), .valid_in_30(valid_in_862), .pxl_in_30(pxl_in_862), .valid_in_31(valid_in_863), .pxl_in_31(pxl_in_863), .valid_in_32(valid_in_864), .pxl_in_32(pxl_in_864), .pxl_out(pxl_out_27), .valid_out(valid_out_27) );

add_32layers#(D, DATA_WIDTH) x28(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_865), .pxl_in_1(pxl_in_865), .valid_in_2(valid_in_866), .pxl_in_2(pxl_in_866), .valid_in_3(valid_in_867), .pxl_in_3(pxl_in_867), .valid_in_4(valid_in_868), .pxl_in_4(pxl_in_868), .valid_in_5(valid_in_869), .pxl_in_5(pxl_in_869), .valid_in_6(valid_in_870), .pxl_in_6(pxl_in_870), .valid_in_7(valid_in_871), .pxl_in_7(pxl_in_871), .valid_in_8(valid_in_872), .pxl_in_8(pxl_in_872), .valid_in_9(valid_in_873), .pxl_in_9(pxl_in_873), .valid_in_10(valid_in_874), .pxl_in_10(pxl_in_874), .valid_in_11(valid_in_875), .pxl_in_11(pxl_in_875), .valid_in_12(valid_in_876), .pxl_in_12(pxl_in_876), .valid_in_13(valid_in_877), .pxl_in_13(pxl_in_877), .valid_in_14(valid_in_878), .pxl_in_14(pxl_in_878), .valid_in_15(valid_in_879), .pxl_in_15(pxl_in_879), .valid_in_16(valid_in_880), .pxl_in_16(pxl_in_880), .valid_in_17(valid_in_881), .pxl_in_17(pxl_in_881), .valid_in_18(valid_in_882), .pxl_in_18(pxl_in_882), .valid_in_19(valid_in_883), .pxl_in_19(pxl_in_883), .valid_in_20(valid_in_884), .pxl_in_20(pxl_in_884), .valid_in_21(valid_in_885), .pxl_in_21(pxl_in_885), .valid_in_22(valid_in_886), .pxl_in_22(pxl_in_886), .valid_in_23(valid_in_887), .pxl_in_23(pxl_in_887), .valid_in_24(valid_in_888), .pxl_in_24(pxl_in_888), .valid_in_25(valid_in_889), .pxl_in_25(pxl_in_889), .valid_in_26(valid_in_890), .pxl_in_26(pxl_in_890), .valid_in_27(valid_in_891), .pxl_in_27(pxl_in_891), .valid_in_28(valid_in_892), .pxl_in_28(pxl_in_892), .valid_in_29(valid_in_893), .pxl_in_29(pxl_in_893), .valid_in_30(valid_in_894), .pxl_in_30(pxl_in_894), .valid_in_31(valid_in_895), .pxl_in_31(pxl_in_895), .valid_in_32(valid_in_896), .pxl_in_32(pxl_in_896), .pxl_out(pxl_out_28), .valid_out(valid_out_28) );

add_32layers#(D, DATA_WIDTH) x29(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_897), .pxl_in_1(pxl_in_897), .valid_in_2(valid_in_898), .pxl_in_2(pxl_in_898), .valid_in_3(valid_in_899), .pxl_in_3(pxl_in_899), .valid_in_4(valid_in_900), .pxl_in_4(pxl_in_900), .valid_in_5(valid_in_901), .pxl_in_5(pxl_in_901), .valid_in_6(valid_in_902), .pxl_in_6(pxl_in_902), .valid_in_7(valid_in_903), .pxl_in_7(pxl_in_903), .valid_in_8(valid_in_904), .pxl_in_8(pxl_in_904), .valid_in_9(valid_in_905), .pxl_in_9(pxl_in_905), .valid_in_10(valid_in_906), .pxl_in_10(pxl_in_906), .valid_in_11(valid_in_907), .pxl_in_11(pxl_in_907), .valid_in_12(valid_in_908), .pxl_in_12(pxl_in_908), .valid_in_13(valid_in_909), .pxl_in_13(pxl_in_909), .valid_in_14(valid_in_910), .pxl_in_14(pxl_in_910), .valid_in_15(valid_in_911), .pxl_in_15(pxl_in_911), .valid_in_16(valid_in_912), .pxl_in_16(pxl_in_912), .valid_in_17(valid_in_913), .pxl_in_17(pxl_in_913), .valid_in_18(valid_in_914), .pxl_in_18(pxl_in_914), .valid_in_19(valid_in_915), .pxl_in_19(pxl_in_915), .valid_in_20(valid_in_916), .pxl_in_20(pxl_in_916), .valid_in_21(valid_in_917), .pxl_in_21(pxl_in_917), .valid_in_22(valid_in_918), .pxl_in_22(pxl_in_918), .valid_in_23(valid_in_919), .pxl_in_23(pxl_in_919), .valid_in_24(valid_in_920), .pxl_in_24(pxl_in_920), .valid_in_25(valid_in_921), .pxl_in_25(pxl_in_921), .valid_in_26(valid_in_922), .pxl_in_26(pxl_in_922), .valid_in_27(valid_in_923), .pxl_in_27(pxl_in_923), .valid_in_28(valid_in_924), .pxl_in_28(pxl_in_924), .valid_in_29(valid_in_925), .pxl_in_29(pxl_in_925), .valid_in_30(valid_in_926), .pxl_in_30(pxl_in_926), .valid_in_31(valid_in_927), .pxl_in_31(pxl_in_927), .valid_in_32(valid_in_928), .pxl_in_32(pxl_in_928), .pxl_out(pxl_out_29), .valid_out(valid_out_29) );

add_32layers#(D, DATA_WIDTH) x30(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_929), .pxl_in_1(pxl_in_929), .valid_in_2(valid_in_930), .pxl_in_2(pxl_in_930), .valid_in_3(valid_in_931), .pxl_in_3(pxl_in_931), .valid_in_4(valid_in_932), .pxl_in_4(pxl_in_932), .valid_in_5(valid_in_933), .pxl_in_5(pxl_in_933), .valid_in_6(valid_in_934), .pxl_in_6(pxl_in_934), .valid_in_7(valid_in_935), .pxl_in_7(pxl_in_935), .valid_in_8(valid_in_936), .pxl_in_8(pxl_in_936), .valid_in_9(valid_in_937), .pxl_in_9(pxl_in_937), .valid_in_10(valid_in_938), .pxl_in_10(pxl_in_938), .valid_in_11(valid_in_939), .pxl_in_11(pxl_in_939), .valid_in_12(valid_in_940), .pxl_in_12(pxl_in_940), .valid_in_13(valid_in_941), .pxl_in_13(pxl_in_941), .valid_in_14(valid_in_942), .pxl_in_14(pxl_in_942), .valid_in_15(valid_in_943), .pxl_in_15(pxl_in_943), .valid_in_16(valid_in_944), .pxl_in_16(pxl_in_944), .valid_in_17(valid_in_945), .pxl_in_17(pxl_in_945), .valid_in_18(valid_in_946), .pxl_in_18(pxl_in_946), .valid_in_19(valid_in_947), .pxl_in_19(pxl_in_947), .valid_in_20(valid_in_948), .pxl_in_20(pxl_in_948), .valid_in_21(valid_in_949), .pxl_in_21(pxl_in_949), .valid_in_22(valid_in_950), .pxl_in_22(pxl_in_950), .valid_in_23(valid_in_951), .pxl_in_23(pxl_in_951), .valid_in_24(valid_in_952), .pxl_in_24(pxl_in_952), .valid_in_25(valid_in_953), .pxl_in_25(pxl_in_953), .valid_in_26(valid_in_954), .pxl_in_26(pxl_in_954), .valid_in_27(valid_in_955), .pxl_in_27(pxl_in_955), .valid_in_28(valid_in_956), .pxl_in_28(pxl_in_956), .valid_in_29(valid_in_957), .pxl_in_29(pxl_in_957), .valid_in_30(valid_in_958), .pxl_in_30(pxl_in_958), .valid_in_31(valid_in_959), .pxl_in_31(pxl_in_959), .valid_in_32(valid_in_960), .pxl_in_32(pxl_in_960), .pxl_out(pxl_out_30), .valid_out(valid_out_30) );

add_32layers#(D, DATA_WIDTH) x31(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_961), .pxl_in_1(pxl_in_961), .valid_in_2(valid_in_962), .pxl_in_2(pxl_in_962), .valid_in_3(valid_in_963), .pxl_in_3(pxl_in_963), .valid_in_4(valid_in_964), .pxl_in_4(pxl_in_964), .valid_in_5(valid_in_965), .pxl_in_5(pxl_in_965), .valid_in_6(valid_in_966), .pxl_in_6(pxl_in_966), .valid_in_7(valid_in_967), .pxl_in_7(pxl_in_967), .valid_in_8(valid_in_968), .pxl_in_8(pxl_in_968), .valid_in_9(valid_in_969), .pxl_in_9(pxl_in_969), .valid_in_10(valid_in_970), .pxl_in_10(pxl_in_970), .valid_in_11(valid_in_971), .pxl_in_11(pxl_in_971), .valid_in_12(valid_in_972), .pxl_in_12(pxl_in_972), .valid_in_13(valid_in_973), .pxl_in_13(pxl_in_973), .valid_in_14(valid_in_974), .pxl_in_14(pxl_in_974), .valid_in_15(valid_in_975), .pxl_in_15(pxl_in_975), .valid_in_16(valid_in_976), .pxl_in_16(pxl_in_976), .valid_in_17(valid_in_977), .pxl_in_17(pxl_in_977), .valid_in_18(valid_in_978), .pxl_in_18(pxl_in_978), .valid_in_19(valid_in_979), .pxl_in_19(pxl_in_979), .valid_in_20(valid_in_980), .pxl_in_20(pxl_in_980), .valid_in_21(valid_in_981), .pxl_in_21(pxl_in_981), .valid_in_22(valid_in_982), .pxl_in_22(pxl_in_982), .valid_in_23(valid_in_983), .pxl_in_23(pxl_in_983), .valid_in_24(valid_in_984), .pxl_in_24(pxl_in_984), .valid_in_25(valid_in_985), .pxl_in_25(pxl_in_985), .valid_in_26(valid_in_986), .pxl_in_26(pxl_in_986), .valid_in_27(valid_in_987), .pxl_in_27(pxl_in_987), .valid_in_28(valid_in_988), .pxl_in_28(pxl_in_988), .valid_in_29(valid_in_989), .pxl_in_29(pxl_in_989), .valid_in_30(valid_in_990), .pxl_in_30(pxl_in_990), .valid_in_31(valid_in_991), .pxl_in_31(pxl_in_991), .valid_in_32(valid_in_992), .pxl_in_32(pxl_in_992), .pxl_out(pxl_out_31), .valid_out(valid_out_31) );

add_32layers#(D, DATA_WIDTH) x32(.clk(clk), .reset(reset), 
.valid_in_1(valid_in_993), .pxl_in_1(pxl_in_993), .valid_in_2(valid_in_994), .pxl_in_2(pxl_in_994), .valid_in_3(valid_in_995), .pxl_in_3(pxl_in_995), .valid_in_4(valid_in_996), .pxl_in_4(pxl_in_996), .valid_in_5(valid_in_997), .pxl_in_5(pxl_in_997), .valid_in_6(valid_in_998), .pxl_in_6(pxl_in_998), .valid_in_7(valid_in_999), .pxl_in_7(pxl_in_999), .valid_in_8(valid_in_1000), .pxl_in_8(pxl_in_1000), .valid_in_9(valid_in_1001), .pxl_in_9(pxl_in_1001), .valid_in_10(valid_in_1002), .pxl_in_10(pxl_in_1002), .valid_in_11(valid_in_1003), .pxl_in_11(pxl_in_1003), .valid_in_12(valid_in_1004), .pxl_in_12(pxl_in_1004), .valid_in_13(valid_in_1005), .pxl_in_13(pxl_in_1005), .valid_in_14(valid_in_1006), .pxl_in_14(pxl_in_1006), .valid_in_15(valid_in_1007), .pxl_in_15(pxl_in_1007), .valid_in_16(valid_in_1008), .pxl_in_16(pxl_in_1008), .valid_in_17(valid_in_1009), .pxl_in_17(pxl_in_1009), .valid_in_18(valid_in_1010), .pxl_in_18(pxl_in_1010), .valid_in_19(valid_in_1011), .pxl_in_19(pxl_in_1011), .valid_in_20(valid_in_1012), .pxl_in_20(pxl_in_1012), .valid_in_21(valid_in_1013), .pxl_in_21(pxl_in_1013), .valid_in_22(valid_in_1014), .pxl_in_22(pxl_in_1014), .valid_in_23(valid_in_1015), .pxl_in_23(pxl_in_1015), .valid_in_24(valid_in_1016), .pxl_in_24(pxl_in_1016), .valid_in_25(valid_in_1017), .pxl_in_25(pxl_in_1017), .valid_in_26(valid_in_1018), .pxl_in_26(pxl_in_1018), .valid_in_27(valid_in_1019), .pxl_in_27(pxl_in_1019), .valid_in_28(valid_in_1020), .pxl_in_28(pxl_in_1020), .valid_in_29(valid_in_1021), .pxl_in_29(pxl_in_1021), .valid_in_30(valid_in_1022), .pxl_in_30(pxl_in_1022), .valid_in_31(valid_in_1023), .pxl_in_31(pxl_in_1023), .valid_in_32(valid_in_1024), .pxl_in_32(pxl_in_1024), .pxl_out(pxl_out_32), .valid_out(valid_out_32) );


endmodule